//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef struct {
  string SEED;         // Input SEED
  string MSG;         // Input MSG
  string expected_SIG;  // Expected Signature
  string expected_PK;  // Expected Signature
} keygen_signing_kat_t;

class ML_DSA_keygen_signing_KATs_sequence extends mldsa_bench_sequence_base;

  `uvm_object_utils(ML_DSA_keygen_signing_KATs_sequence);

    
    // KAT arrays
  keygen_signing_kat_t keygen_signing_kats[];
  bit [31:0] kat_MSG [];
  bit [31:0] kat_SEED [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    keygen_signing_kats = new[3];
    kat_SEED = new[8];
    kat_MSG = new[16];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // signing KATs
    keygen_signing_kats[1].MSG = "fc2925c28f99410b1f0185546e7219797299369d27c6ab2d00adc627ba5564816fd47ef3175a769ae51fd160d23e458403e27cd6d16678ca6367a098d62e6610";
    keygen_signing_kats[1].SEED = "1beb2f2b7967afcf76cbfdead98ccf7637b4aef67aeaf2b263a324bb0885ed3e";
    keygen_signing_kats[1].expected_SIG = "85BC06C0229185010B1E23D65F9F974FFA0E86E6DED4CCEA6965313028757A7C4B10CE05BE1A3C317BE542D87EDDB3FEB57B785F28071772E2FFC49D151F5E5506C0B21FC934B6ECDE9026E344F18B21945DF950464725B94F5A8833B6185CAD50814B5CD16A9CBF44297426FBDAB19A9254E78D0944B479E7FE6FBAC48DFACD8A15DE627A60BA177A5A0445F84200B28330DAE2BDC30A67CCEC75A53BB2724BA2F3CC0CAE65FD48FD90E02524D3657441D376EF59346E64C2B26556C782A12E9ABE697BF58A70C3DA3C3C79FFCDC6B290F5D1CC660989CBEBDAD2094E96508EB9DAAB000F136BC370CF64CA556583082C9C953495C1FBCCCF6A209D546CE998425E0E17D81018153FEBFDD73D870D632D1CAEF5415B8B00E1B752432069139F514586E1ED7E55E695AC725B770854FA78AC27D75809D7B85D615D7092B2E609A9C8A9347623E3DE0CDB4AA9E782A4367EC1799B02106707A44C60535ECC6A7C4F59D1406900C3C566174D647F249C4FC2C4358EC5D0824030808F77CBBA8743B4410432BF93B9771BF5C92B522AC368C58734C0ACE50C3295E8F338CB92E9BDA9D4976BA2C60F3975DD074A9E8885A0069E92F839A26BCD38E639A79369F6FEE8E1A9CB0B2BEF03E196EEC6BA0838336AC40BA11917AABCD71CE8F00437343483FF27D9BBF2328449EAC9EB1672E750A79E3CB8C4BFEAEB1B106167FA56A8EC9F506ADF953D1E2221487F190FF6121541C3C6D3867B18DB63FCFDC279F2983030DEA61FCE0DC8F9BD0F8E2888ABA0E84AC27975B637B1B5DE12FD8CA9EA1E64CA16D845CAB2280BB94BFA0BB4F39586CA303565104BBE46A7F6CD3AC14865F5CC06894B2D11D26B7EFB845E9B9E98D3A6C7EABBFB03A66D7F5E7C7B210B8F240ECB1B62CFD4949C5352099FEFD45076B9636B89027F5596884C2F09A0851060146F575F4841701507F6660A4209263B0AEF5F8255E98E34BD7687D5D554CF68C6C267B1B1F10AF6ED940FBC5993B924FE925A3C43E2972BC9D00A4F13716B6822B34E165814C1C98FE7B34ADE716B21B326C2C0BC13CB86B9551D228E1A7BC9AC95BDE1FE822805C9FDF6332AAA10838972F87CAB9D160DF4C1E7EEA533C33646BDC5EB46234837CC5D46D6957E1F8BEDF493DBBA305B96E46D3FF39CE38FC2C013C5D5C4946A8A414F4C68BED207524673DF40C449D087A1DCA3D1A4BF0F2F0FD139528A95E2BD33072D125E31A99A17A1977B8BD58B652AE870D6CF743A52DC343F9D4EEAA10EBE2FE1EC57A8AE33A2050A40697B6D41E881471A8E720E9E39E71DD72335A6AFBE743437061A522B9B129DA4B74033356D0E1A9591EE5EB09E11FDCCD4E422CC6759B8DDF118A82FDDC975C7AAD69238255B1713D6B6901FA5E6411956038D831A077A8D90556C9F6CF48098F9BDB838AC7216DEAC2A84453B12D26B68C20B8EBC8C09EE4FAA40DA772D67FA8B474F9F3873DB8CE4EA74B72800128D94B5DC91AECF35EE24DA495459E2844AACAD6EA69015B7DEB23F06368260329CAC40AB498217BBBDD89115057EE95CC6BE72AED4D7456D897C7DFA55609FC4EAA162873E307FF1E9D202373D8AEB16CCDD45CD6BCD3D97E433B5912B2CBDA5D3DB0B2CC103FE7013128CC798B97141EFE1F888149C9F007FD02EF6F8999FB1C1F404793FEB582E94ACCEF2A642528A66A1DFF389E2360035EF98553A2F09B19911200B05DD8D781D9BE9D8191493678383C52519A5F98BF63A9E834690729BB9EB61834AC611A64771C8373AA27B3804B0A561CDC64D9B986AFB50C99B1F1CA07783F06CB8C2CCC88490F6C5862DB10B9D61752B0B03D2D93B0692D5ADB9B3347607FDEF6D2311117D28FEFED7738FEBEAA589C821CB2420DB361AFC5537131BE739DC9B7DA2099AA3DBDF9F04AD245AEE3E065D21848BE6E1E5F87D81D4322BC570264BD477F91FF0599F4219677CD228F87183C5249AEA2FC7FD1239170810CD839E4B8158B6595A73A96EF8B9E065FF5362ACF2AB0DDA13B0B9AD43D88986C664E76849F98C478E1D52A1FE4541075CD4229CB68A4385618DDC67FF635E477F409811790FEB183806FCF63216F36B79AB140FD39764E15B5C22B7D22C34D6440F4EB10BCD72E4F1BCB0AC98BF060FF857AD1CAB1539E51443B214E6C6BE287A5651C6A33A7CF8BC3E5CC6C09C240762EB2F0B25C80E6BA866F6B93696113C9F43ED4709BD7221628090D19BD575BA654F291A83053B94B47DF9497719F91296D5E08BFA63212ABD24E85556663A35890D21A97CB8A1A8E0DC45653093A058B2DAD1A0D1EDAE2F43CED4B84AE0206A77B6B35150F544E166CB30E47BD594C452349CCE2F71327849E334146CC5662F5D057E689F7AEA1FD2B1BB0F45BC04CEB801514F3C930E44EE4EE93ACED39917695546EFD5D78C090EF1C2C1272A87ADC3646881EAE493CABE4E364053AFCB22A621BAB938F1B2FE8393E84B5D2E113B51FDF720084E4E82EBDFB894D52C264D85AF5365237FDF20A9B4DD13A384AEB1AFE877781FC1B62D99878CCAF5F4B797C96056AAA11613719F60E56BF3AF4C0735A3E1B5F691129959A0ED13D627298EB461F7EC70AE9B191F2B507415119BBCC4DAA8024985A7D7AE424DA992A2587D109281B183DA90813F287406521565E26B2645009870DE574A8D0AD0DC73DA19F26AA85DFECB4792254E3EF5BD65ED32B8A81C152589F61A3E63E2B7BD46B490CCBBF17216697D5D6D87EE32545F900F5983CF3226DD997216897D556DAAD0D1FDF61D78378B5E4420E10F4D5CDD83B2FDE4BB24C8D8119F48A912E8BAC57D628B0ECA5F7C86A06925777834141D2F7B5B317C9907947166963B77059B7AEA5680FAB0F0DEB76AEF53489019614B7293AF592FD485D61DF6C99F5F7320D56554060053BDAAA982E89FB39DB5FA03C1BCBF93C2BE56FA310A15D85DEE86613DD5936D9020435D81795FBB811FE88D85D369B2083D24933443C0CB710CE29F50FD52A7E1209AEC6CB42EA18298DFF910A216BE1741AB1E985304CD63F1C2F3B3EB578C34BE5A5845AB38E91C83B68F9DE9A5D644652D60821A77076EC17A0A1AA776498DD51B95811CE82B2963D379890909E39E4C1925696449BF1365A8DBBCA21D791DD64C45633A596D8B6B926C4015F114D646C3304337560440611F7B0F87BCC4EB659F3667C9D3258EAF4EE3096EDAC3BDE0A2DF61624A318FBBBF1FC42E2E70017E83CFB812E374F1156B10F4FB6CCCB2E8BA6AA0B7BCC268F3044014C1EC56CF3EE0C8641298112F9004723E5847A4545FD34B9FFCB4124029140D352DB3A1E537A93E70C9E93A47B80979E1B8FA48CF44EB6ED479DF6ABE93BFA0B7D3B47E129AA9890302FFD5955395DD1D9483A627F530E8EC59E1CBE0542A3BB93DBEB737392FA9444C760CAE232C35D16AC8AEF4DE3DC5E55B7633DDFE1C0978E8E5D2515518EC5630F0A9F671F13790283B6159549622E1766D641E609CA26C593999A7ADFA8214D2351E059450094C54DE934A28E0D51F59FFA18CFAAACA94B5A1B9DE5539F49F9F0A790ABF8C3146A1B87038045C7F4A81694B7442420D9F6456E820FE081594071831367F58C1879E57B44F31E74982D66282876AA3C9693BAC0B81406A24E6DD94F3076D89F78407B7666A7509A06F89152D0B781AB6654BE96908E3B667B88A8F138BC5DB62C86E287215D0F5D8E9D4CE3FF8637F86EC85E3C73A9BEC26069B5B769CC446F87110BBE0BCB1B53BDB7DC605666AD9B23B23BA3F77FEF401AA108DCD298C751C6D901B96ED34178CE181E3A09BD1E98F97BC8EB21818D790E851C2CD9602A45AD63CDE41354DD9AC3BAFC5ADD87919E7CBC82D589D26DC0381334C104CB9B9983B6C2E10378AC1310F5C412414D5A8435E2C7DAF6C27DEFFBB1AED3CF135429DCDC0F0F5A9623EFF31F7EE4FE790CC46F9716DA34A15AD2162AC69C216F0F3715EBFF25A6C71839E54E14263CE2C7D8F6AFD1C6B7EC772E0C0EC395DB3C905D5BB5D8E1D3566C7B2410247DF8E730530EB9B9E924599D70A3E9A6C973BB2861355822EA7CA328468EF097A5A3C068390E17B8078A4DA364980DDB80A12C2FB973375333E2CBA83FFB331614410CD8B9554AB90EA4598FBBC71122FD7563C5CD69C3511F20579EE772671CAF34298F6369D8F2B5DE0711F4E145BFEB75E8767D48D43643695D36336C5276A9A5F629B7D6568FADF26327A69E95FF267278043DD9CA0A4206BF9E844ABA3AEB36AE12233FD8CEF1D24CC3B96AD5EF046F1975D7298D99A76BD949B4534B93C59CA7B9E5589EACD6173EA46A9F7FA0DC6588EC4D4073734D0816C6CE1260F04A67206A997F9CF4EF23848CF247DD9C2908FE15B1CF1904A4007B765DBB81F2FB1022AFE5C93A612DD70A7490BFC7470109AE1AA63CA69D1CCDE9086E9032A71A4AE9A3A8574B67029D830FD641392CF60E650515D2AF8DEF25D3F0C070BBBC7C16F94B214F32A7668951CE5BB795FB66C3E65053BBDE5CA90FA17FC02EE42DA713E94085AF9C742FB72041B1710C91B570A7060EA322C6A39CFEE0850E00F019945F41A290E3697CC8CD8C9C85A7E3ABA7563625BBBC2B3A8D344AE187701BE4D38AA5BA1A5B7011C250EADE01E2A12E4E75246D2459C06377C1427DB30563B47102393625729C3E12788683483962E8E6C6B4F5923D360F67BA39689DB6FE52D4E7CFEB286D6145C3700573F62470436F5A75B20D0641EF8456B670DBF8BF0C022E76C78664304C2589DD8F158A32B57B9122C60D0680AB386B3732F430B1C9D18641232FB322C4676EECD203790099E2A78640276C37476A32F72AC89D9CEFA40D438BAFA9C960491DF1CA4C0574B28EEBD15DE1076DAE402BE4C5AD88F480923618065C6B00781B79C149BB7CAC9263016F8B8502F6305581C94C693D655E84C9BADC91E7EAB1D1E987AA9C4781CD1E2D2DB1FEF265180B322CB21E62B915C05CBAB0AA876F3AB2F44B93DBAF59DEE23338224F1F62A0397EA6034AE04F0C6D5D6BE4465B8FA0683695B5F2DC76080F9A8F91BB8B4D4F739A5615DEBB33593750877AF3F52D80FC24C9D79957AA868291C91E77660EE41F3E7045AA53BCF5275BC5D9C821FA35B8B05CC8FED3212514338E56B07A476E4683810F7D5A35FFCA3A706EA218A40241C395966F99A8C1DDE202CA97E11698A0971401576264A5836D2ECC827FD4495F5667318FB73BFFCFA330A9524FCD20478B0B494CD9C18C6CA5C8EE9E5AF9DC90E25C3304F543E6DF69FE3FC3F19B3F520D19EC2A9FE49FD405244763C8F94E6DB9E6BF9C2A614A219A9362AD2DA32A998C2C9A2FB0B6BD1C0FF892E0EE163C33C9F4B7E6ED91940068571678D714BFEB48388AE29C66BEE27D633B50D26C571FE969A25BB755CA44EEBE68E01BD1FA9A175A5D2C1E0838719C2A7468AC9051DCA0569F193549443D77E57DD83C66BC5753E71E4E49853CB6BBFEDB61F7F0645B4E0A71F16DDECC2C371CAB4C2DA3A61BF27FF547FFC512B65E7F7F0285C9EC7806D615C8E0C3ACA1B762DA6D04AD99726A80213E0B3185C0FD09697B457CC1C673E87ED68FD9F94B58AD1DBF680BADC2C4ACFD970DE2C72FCD45E2CC92ED398E43724F55AF0F88334E849F8B0070AA4410A00A511F114C3AF05EEE66C6CC6282CB6C631236C1BF429175F632972AECCCAF29DA563610C8EF04CAB5463F32A8FAFBBF5FD81F399F684EA46A0451B16CDE4D101040D36C891723EAD87C8A9B1245459A4311BBBA2464F823ED60FE42EEE23481A565E15D5DBAC132808500AF67FF7A93998EFD772D231098AF4AEF6E9FAC876EB89CDA56071B1DFA5FB3EB16C97358997FE22597A35931DDC4C3604668A7A3333B24B7CE50BC3B2A073B3AB537D0A749260998263477A1B94014FABD8EC14B55589038AAC001C1A4C395EC4725CEA619A95D93C4DCCF61FE9FDC8714B112C31592A8A226E364B13FBABDED4C2952D93DA4A50F7FB3747829F613F3C31262F0DBCDCF14F8B9A5E82D989C20AB3590E88B4B6D6AA6758D736336C6C1C9AB627EA2E97250708ABCED1D2ECA7E16B8AB1D159363EB0091E1C4779F6580AD7FE78AB31CA96A822ED0E5F3469261C96391A99BFAF36CF725F24F815405EC1BC1C2DC7CAE945DF5C4F54EE523307DFC57E89B700383B3164A1582BD61F954182E09BE4ED83123346E0CC969A90E7F76B9CFB9C9FE55D6D0B639F5948DC98C389DD3E00C68FEC356D2BADDFAB03BC85181293467EF674FE919A8C788B1AAE1A71FCAF47198186692FE848C77FA47944B33BEEDE85A9D2C51CD9621A49EFE79660277F207EDAABE36D068D7BE36A0E06999D2F764E891D27010108D64FED39B3D8306AD16A62CF45D8AC7BD02E9EB1A05E0869ADB8E3C69CE295CD1642959AA9B2C2D72024263045676A77949FCACBFE031B2BC8CACBF80BBCF70F5E7B8E9CACB3F52058595A5F858DC2F8FF05137D9FBAE9FD11263150607A9BC8F0F50000000000000000000007141B1E2630374100";
    keygen_signing_kats[1].expected_PK = "3406C20EA187919F41CDDBF27F9C50A52B7EEED2870011EFF9EE10E8F69E0A39C794F3F7066E3CD63130D93950D0161F14CBA67DAE6D13A7DC8D9F439A6C626AD4005F3A48BA2E531C42E444E0C076496BC07DD0644D7096082258AA0D37F3D3D0D587E0064CDB9A505965691E27D295802D856B3295D4EA6562FB3247E343B1AE264E88A02B2777F92B64686F3F10C833A87FB693BA1F4DBE1812BEF2028BD37625D70CA9667320B8FBFB8C390BDD887A318E7AE9326BE4B457A612932C934E118ABC31A9C79D585AA4128E3559FF8790B96952C372697E96FAFF01E55168EC199E92A1360C3AC2196236561DC697A0599C072AEFD6A2683ABDC3C11557EB44B936465E15994D14C9B3F0E84EE72949CCFB9531F8CB75D79C9C2E68A1ACDB92C58A9C19241388C054345CE46CFC8AC2F1FF328639D09C071EB9E920F697943145B8FF45EDFBD8F5135929ED18091055CEE48E4776E87BBD62595E21990E72E5C09F48EB6F311773E523D395374AB1E0CC3D5B55F7EE22D2B189A882939CFE85694682685368E272DA8EAD2CFB972E4616FCD8143782C5C3A97F51CEFAC81387700C74D5D2E5B92CF762A1F327841AA117694ABA918FA29300C27DF3029EECC775EB2EA2E9EFA882A0EBA9E82C588DDF09FD4620E084756F5069BE893CFA1D8E0EC69962774E70D41F46F25F291C091BBAA447ACD24BDF5E7F0D6C50BCE69B79F51A4CA8FDD8343C49DE55EB3441E042404CB992803C2494D5512AA67A4BBBBBE765AD543C709A07EA71083EC4007E4828C58187C5FDCE680B34C902BD902A85E38C674B07D13E5BFC15CBD547867A3CC9A00D0DFC5219CBF4E82E7010B009493EE5672BE249DEBF2F4E91B5469F7CAAA5D5C69A080C8EF8394F06B8AC95FC8489A0A7BB21CAD3548BA524B609EEF7CE7C20DAB6C5B54B58307B416C3DB4D653A1446F25A8874A7B8B0AC6C2DBD175726849265103D455B1895213BA6C3D177CCD788145EAC23A65AFEF9CD75B0C2F0297420CDA46AAFCAAB92EE9955948A741BC3F60AD609A53BE44624520252957B2BA03113F6FEEFB690D0A7F5952FBB470F3F9075CF9EF0541A9B6BAA9DA6795BEDD8F41A27DF7F6C5855030354138E2077B4B2DDC570FDF0186DF23F077E1CF6EEF833D0E4CDA82709B69F9AC52E4D9254A7D0DDED46D64EF083C3585FA3A5B25D0323FDF17EABCBEEB64BA8513010494DF411045DCD48B1565697B0DD507450866E582BAE23C15010B6088806C254E6D81DFA7922F189F3A7559792F198A96916F96F78DB378541D02621D0EBB78C72D2A360E47EF09DDFBE1B2EC24C99C692E087D84C0BBBD8FF02275B51813624E97448C5FD294A2740D0775060A8F785630402DE3CE4357A655CB6DF2C534FEB3DAED1E1FF7C6161A0B0718DF0C2B3C228BB69D0D8828B876114B95621EDA905766E877DCE20756525A4C31FD84963974D984043B5A4CABFAF21297390A09FB6EC15867734065C7EF6B18AF9FB3596919820D21B766F5F2154E8BD3C74FD711C2F80F90431A44AE34997A9085765636D27CA3C3A7CABA01902D7554B0FC97180BF6547E97CBDD5E094CFF25206BAB14BF30C41EA76268996D4F011946387657B61E8715DC097DCDADE05A72712179F0A110E4203086C409090371BD175CCEC01DC33A7F4F20EF3448A1757E0C560BCD7747E6177346A8B8BB8F9FA7D04BE2D897BD3D5B5FE1231059BA5BFE40180A7F3ECECE7885B09970B692548C3D065BA17522151E0EEB32F3664C67D5164F92B48F3E167D71E11F3A822A2585BBE6395A9DD827933C31B7E43188830E5CF60381D6CC58DAB278AA0A5192F7CA4497704BF951000E3E786AD4AA651CD9E1650D0BBEE5B163287B44C1A918F6AE43C14E97A10E92F3F5F8596A97CC54094BFD618D72C433E4A7BC1ABBEA4406E5C5C8EF3FEC6F750CAF9654295FD26AFD89BE26B000B33C1F70DB955628AC16C0A25216942460A61A6807131EA5396ADE6716993F6D4D178B1E604DD078F2B488F784921467C3F93A4FFD2B9936F1C913F48B51EA64B64371EBC7B0F8A0ECA57FD0CCD614A130CBE5B9B2736CE5EA9652523AA2033DFF532F9FB94685456DB9C044C9DBFAED8B74CC7DED328737ED6D7CA13E55397699C8E0DE5DD7CA508EA4659C21A07968697BA3CCC7C9330CB7F8B95E7353D2B3374771709F364D82F3190134A27CD2A34D61869962F2403CE1F3218D9DA220B540F907E3AA578DFB60777A3109339CDB7304360E2754B3D07E132946C9DD795688A0704C75B10BFA36BC1306706353A1FD0BE5AE1560B7903FD411E49620D54DCC194D6E240FC87712C005D928B7A07C4F3337050D6060BA51EEC1D6FE0D7D73B39547E5F9331A6ADB3202EB2EF327F69C4A4AF35ABDE056475F4A4DF8728999D4D4BAA1650967269063285456D4CC8CE8C1F5B9E29E5305E387D34FB7259521E620D68DAB8532CFBF1021BBC8179F9225F38A0F04F19316F388DA2C4F6BF1C8F9A6343D890E4E4C71BA1EDB0B6D0B2FCCC559CC20AE06352C75E09A19A109BA1F1DC8D5CECA5D46EADA1AD47BD4F67FFCC40AC66DAF5B4DD15658B618631861EB6564BF13E9CEEB38225715E484983A706020875295D9BB289024EF61D116BFB84D72DD2D0F3C0373CF0605FE838B18E4A5D8DA5BD23D9E6E2B06E7044DB3D0774975FAFA8BFB6DCFDBE95EB5262FF93663A0A6F8A7B53BA1057E611FA1B3A3AF42741F291189CE1E2F628EDC1738767B0FEE93E66BD29FEB1C7CD9CE2D516CD9488FF33E9CE52198B05E2CD25020B37BA092F962B911864AEB5EE5E0037D9A5FB521EF99A1120B9A9F68A513C02E72794250333B68CC3A0AB9E473653D015CCAEA2B102B332B3B4BB95898440D6D290E73FF8F80EB40C2DCFCE9EBF64C574EFB9A1C3BBBC5AFA4D9F05F36BA6B44E66AF4959B79D706612CA98E689C56DB11AF684A004034FCFBD106BA1CA09D97D51BF20E2058FEE0E1A69B4A60B9834539AA94BA63EE1402CCF0D19B280109DC296CC2C40CF8441BE76C7DD2D17F3DE72B11C4AB7883FF352AC5EE4630D37BCD8D92291913F4B81021A094FE3DEF52824068C5FDCDE8EF26976B29DFAF51612837768A69CB3D06ACB1FFAA0B6F5FA0C5AE618D2156AB91F72697323A9D8BD3FE24A2B884B635CF933D2F80EB0DD48580ED87A30934AB5E7A5899299D366C09E7E3215935492E9356E3673E4DE1B29625FAD193BB53C0BC88BA55788A9970CC007288852661DCC161580FFFE307BF549F2721090C5B6424E9FE7852B8A76C6B06E9319B41720979D685669E95479467336CD68C06B48A6CB6916BE4D882D0C6371380F97F9AAE546AE520D843514E315146C7599DB5DF4D4BAA79EEF3EAF8C38EEA0DA201DDC5A954387C372FA1686F52C8F5CEBB9D54FF879D7339B5DE8BED40889DB44FBD9302BE8F0C20CB945389FE9B56770EE176D2999A9035DB69D9D13EA4E6F9CDCDFF55A5B6945604562915EC7C81D5D2B49E5B1750B01051E7532B8D644CADD714512948AA7F2D88CC5F154989A7D4221C67DB0852C02F6EC9A1EFC7CEAD302D871600C57CDD3EF134DF2EC0070EC7F8D1A80919045D1E630B426A941E15A0E1D6E258F47E2ABDCB9CA791F99885867CE36B6A49DA864A85A0C82B97959B";

    keygen_signing_kats[0].MSG = "ca393154ce0e065793750cbb96156c74eb704ed0f2ac97c1131f250f550e1efab980c2cb146960dd7c0b562a1f412c6b2cbd203e1f048c73376590bd39d7a969";
    keygen_signing_kats[0].SEED = "2e693a2372d55bf2e3793a2d54a7c9dd70b92c0c2f78bc56450ce98816c5f730";
    keygen_signing_kats[0].expected_SIG = "8A659F891085C42893C7523700527092698C1C191B0F187A493139A48BAF373B92B6E6D9D507A0BC0F9CA86226FE5589EA760E99F2D4E22378E4CA968A3E945F1D7F36F97F7C11CFA5CD67D63EFDFAE7DF68DCB8A3D6975673EBCED7D8ADBEE342F7B8E6F32E6420B520FD284F72DF044D322B15079150E6BC6FCBDD3EB6FB175238E3306069B4EB7EE239FFBAEDA41C704BC3F38280DFBC2EC22DC806357E4282F41D3C63FC9F6B3B0A02AA0BA960A45066424A59DE99D43934B48BBC28C8E30066214A1E13A967D5A5CFA25811C013D85BE5BD1490C44F2ED16D7594011AD2BBB4339914E650A604B907D8EAF80FF24A42B0DB618D53C14857344951A653170621A225A06F70D0329C3EA15798A28C1111C2E4902DE9C04C54525254792C5C0DF0668F2DE6F3D77CDA05605A7741A4BDAF5650A76E68BB8BE505CF1B4C18EB3C3820A7A90E69E5D170C87DF46C29F1E024987681A1D36D69ADC6879C0BF785A8139E2A857DD4A76B29963DD28ABFB9415D7010B54A496133E5BCEFBD9504C0A541A3AF30A97337B249F585F604580333D83FD453E109442E1E0E4E37105781F4FDB9590B05890538BB61414C3094E0E110116FBC25088F6E32131FFDF3E9AF8312D603E25B695D8F6D9918DB442BF60F2C4C8F395A7089208D4CC82A99AF093EE32C216BCCC4E799A0FC9A9BBA09FD372FDE10F0C448B4B9DB4631D03D9EBD8BFEF09D686DCA17D1B14459C0190C4CF9EB53F47F4E95768364CEB2A9A36CAB718BC483CBDDA9BF1AF881EA346EEF7BF245E09E08D3F355AFBB0B3F6420C725368E5DB7F6182CAB20C82D1363374FF9E18F444111923E94BCFCD236293F4E47C391184CE4EBCBE1716B1638B879F7D526A12C4990B552344570552E0647602D0BE13F4DFBC87C104D73760EC31EEB9C52AF2BE770D73CC4794A88B61F2619EA0AD19E90BA1BBA75F8892977F3935EB3273AE04038B94AE7C3932E10B4D45E24B5EA4E7F767ECB2E929CD0C48DD5BDEF58646A17A15961FE57E008DC1B5E5331C8D2E3CB3A3EBEDF405476D33A53D707A38E9CF5D9066B84DEB8AE8A75CD776877B5C44A90694A970614E7CA109BCA9B76DA126C402F814B8A2D22CE7C2F5CBDB70C8A0595F922341CF32307E5E69030072F91B32C29D1205F0D585ECD2862389A16ED461E0482F65B3063B093ECF46B603863FFC85800041650143D5871660DBA750F1102BAD4EFEB3DDEA86AC29D0510E00B5A811586102A667B76F997FD6F0A918782327CB374AAE591ABB6175AA15506141E54E622325DD65E4F4C8F69370C6D82F3BD06F80B04DFDEA8D547B1A2AFDE90DF654B37AED1F1DF080B24BAB6C3D337A25720AA73DC3E5CCA88F71078B5D3F2BA1812A593537171691DC313E21E9012ED9DECC6D20416F840E14712D6AFA552022C7B5EC578F42BAB2F77661B2C4754541252251B179FC765DD52A9556C650E795CB153B2BE5BC8AFA721F87BDD996F7A82BCE1955F163B6B951F837E5FFC758FA92AB83D472199DDC8942902713D15F5D1B57EED176AF6366FE11932507221963D8D332911407F04AB610DCF434688976EC347B2B6748515C82329A3A5D31BB3D5A73B0959184B1BA8799ECBBEC94B5B5DE2A794810AAC46D94E2210094ADE4807E9DA3F26327A32E019C52044D80CD2502E67FAAEF5087ABBAF93543BF9DC3D3544163C469952AF12670BB21CD946210E059DE868A52B34BE30BE951DC81092ECD0CC261803E25B7B56F963D58EC92399EC96E095721E2A4B1AE553C37C90CA8EEDB76FFD1CF7F0B7223E6BD68700D2B04626D12EFA1053C65BB14892C623C8872B006F8F654009AF571A6F91D83AC8E6A3260FF78F946A197035BB4AE04DDC9BF783D315EE35ACAD9BEA041E5C631D2C860D4402A865CD3D13E82A0158114B5F51D403A769277C0056C4C645B29177B79394B639074E85918E4D9244EE4C2FA2E1DA05903A516C5054B348FAAD38696DCA8214914241F658A0A659D36A96D96515D055C87B2E628F4FDE39E18C2D0F164DD1893F3E595F11B5463117BE1EB276328DB1073AE17EFF6419652840CF7F99B93703C1FDFD41102B02AA6BEDCFFBEABA28AA3BED6FA8EC790243679E629397E64384493598C433E5A34F1A96EDBB9697094D16F33F1344608E3122361B25EDB34AC763049F5EB9D21028553893659049AC318F6FB55B6FFB13D245F09A413D06C6D9ECE959C2FBA470EDB17A00B9432665A7AA223193075D7CA97B2298437F77F21775F8867270B9829CF8BD7CB76BE6C6E8F1036BDEE6E2DBED599836A43432876B44BE2930741CD934E5D0291A8457BF0A612B99D51D6CF4C412F5A156222AA1548AF136CCE6A57D3BD730D0B0A3410F4303187CC23E6032DDDEF14CC65B45671A8C0EE608881CDCD7F558ABEE9714F25D5C491068E3E278CA01209D96EB6EC8C679B21DA34AA9B494B4A67F2C742AEC06653FC66D4013557AD388E8EF21071FDF117102786D4F2DE16A68BD4380BD18558BB29FCE4FF761DC3D5DCF48289198B1DC586EFFF23FC9A89478217B37FB6F69CEB89EFF9DD0E045CDDC05A6582E277052E51C65C6DC5521E2F59B854694FA985D05E923D14BB7EF6AFE34E63F25DAB21F669AE6C6A9CC70BD8FD72D30C9224D6ADB2F5428193C6190BCF1C073B409B0C35B658ECA358C2B9D24D02E5F5926AD2329829926C3F39B0FD49BBA44A9D3C5966F07B4A06243AF5CA160DEB492E1EA4847FF4FD14CA75B40D125B48ABBFC3E5B764A19A1D491AF110D876FBA529D3B5D3A3E48686AA9AB26947F1FA93D9D40C3DBB36FF652C7A30A3ECC728E94583DFF9AF8A275886214B6AC055F3323B9AB25B3822DD0C2ED64B95E3DFD9E4F50D547BFC790694F38CFEC4146DBD8DFBAA2D78B2B3E11F340ADB8BEDDEDDCED867D584F67B9F3601A62F2660932901393486156B0D61FD6E6B459F5C01A485979797F1635687EF246C960D64C1A248145F5D1658C27D42F0169E71825EF9AD8893673A5D323A05D28E444660ABC4030BEF6C66EFCB057A9EA0684B1B64735728DE008A65E2FA43B84CE5FC39649AD06C92119DDA9C70DBA340FC4C27DACD809637D4FDB0634684C5936B009B5FC3FC7D9B09B29C70ECFF695D885A35C21EBFF236BCDBFED085F7B4E609626221571C8112F03748DD010FC97FADFCADCF825B0472254C026A0C5E83610E870F75988A7148F2BA399E5891164E59740BB41D6E6277C73B1412993F91C3E2DAB02A4F12C427ACAA14B21973C1D442C79D2F038AF9AC48A0D5E12EB82E234615BB8692DFEA8A98D83CA3DD9033D7C48B00A0731EB2DC01377184BE6F2D7DD697D44787C6A6053E6E628437FFA0419A0BEA50FBE52D6089A71B2E82D002EE1FBE6BB3108CE863A08E26890DBB769A417E8926950419D2A952E20AEA560EFD64A525B63E46D2604DBD2CA4EF862BD3096392D5455A21095CA663F886460F592BC75555FE9B13A00A8CFC9D6991488AC59CA87B8A33C472866F821D20F99BD228509F561458CEA2D7EC30048BB547E53DC48F1F976BBB304FBCD3F1DA708941A3B3EC3B7E9992ADF216FE127CD16E5E23B08A7E364704184F659DFBA2719E3C78CBE2F19CD4A84F12D5F60ACDB839DE814C52D30CB8B216A443B2F98225C4E18653CB36CFF848C0E07FD925570040E60B9810BBFA1FF2FC92A0F9EA3E3C74DC443D5363DBC576684182B13D573BEC531151F32F94C1CB54533ACCCDFE86DF79572044054713F3A83275D47B552CC7EEA9501DA6982CB81EDD982CDAE683C10EF122BAD67AA2B69E1BEA2F628880688ACC773ACC727B0B33B190EE05F3BF5523C610CAF7A838A7B9C3F185D44696649D354E1DB65D76832EE32BA1749716BC509AB60688164A030E06B5866968B3CD64E26950B0BC99517219AF04AF5B79EB593B0FE4EB497293A688741027F0725565677ACC6E9432901ECAFA14DD2611144AA5F4F0278DA0F9D7502ACCD271DEA06D6A89C42D473EBB50AB9087202E8ED9E4C1476B48445E3A7A3E022F32A220BF29B5442E41E0106D560EDB47BE768D620B13767EE72E0527D07270D2178608FCDF80284668CE9B74CF63DA78350CE9BC7CCF87B38FDD5C4EEA3CDA098282285D14B74072F07524B0E68EB7E780EC225D6EAECC1DB7610A757508D752E3AD82C5D838B72677FB78EC5D5C0A6010BFACC9AB90CD159280F440E886435FB8A525B8AF97469A8985211A83FEDBA6A06D713868D544F104994EE93EE0A3C42D5106B6765210583AB868BE1A5B9A0269757CAF882A4B3C2D4FCF8DC4F3BDD409684D17235763013D3939FB4BB9197175D6B25A966399FA0BD6486A63E4A20B91B987E955CDE99DED263A9EC0796BF3D14B2DFA3BEBCE7CED3E0953C02A44596B4623FB73F60C6BE64F0DECF9D555CEA95CE07C60AC56CC0C20D9E39AAD4B51D94682C0B09010E9BD1A8D24E1BBCE8FBDDD30980F03D67A6413B95C22EF21B4E889ED43F55D787E2CA0CE1B3E237B46BE54B65CCF93E05CB4D63141BFA54F90CCC5B239417A8AAD7A88FA7CCDE45B26D12A664F49A8154A3965FA8E3CAF276E35B6AF06D8F271CBC18C17253C0A7E21373E7CAE61F6088CDFA4FBB434B206D45A3B937DABC331342D39CEA1FB4C52FEBBA4F89136AEFEF338F021E4AA3E0E028539A5F126EA37A1456655311493CF992ECD7602E150A290EAD12C9041ABC57C13EFB1A3ADC7F3ADC7690C8217B85D2D9D92AF969EEE20960A74759FC0B91503A391A7CD57FFC822CCEB8CD555F27C463F486BA2AA96FB2776EB88714B3225C3690A108D14406D6BD6241EC15CCDDCE4FDEA4032A667641144716BE03D02B52BC002840882B9C377B2BE19CE16A49867CF236ADF14E3401DF348A642548D36E9FA1FE56CD02DDA2CC05A50E4BAB45174A8BBAF0DFD8A2662E96DCE4F823509B2FD9172C85C46F281EB9785D4C9810B7DDBDF984AAF2838D7C854CA47439D4D359A7CCFAD80D3BB18D843818A0F6476162AE74766C55F217E2F62230EF763A34B360C7AA6B3C531D6869800AA8D933B7BB0E63FC942DA2E9B194BC55FA64ADCA4DCA0A58E898C437CA9D1239F50D9CCC834D9DF1E6BCDF8EEA63609AFA46852324B31B96FE4A535083423D59560D1AFD42F3F3C57E98DB0629AAF087283DE6754276173D3BF388702E263022A30A224466433239E6F0FD13570C6B96C491151EF1916EDC7865E2ECDFA2CD5F32332E224757E27C6ECDCA51E34C498D42BF07C3A7A36B24EA3D0BE1D668BF5D011577068C05A8EF206660B3460B252B39F0BE21122CC46541C4F79148D6099F78B2F7D79A2C8E0477DC2D19E0DF277E2504ED60808553640BA21E2427D84CCEDACC2390901D4D263BFA2BFBE18596AD80DC44AF44E7B2D0F41FB9EA0890D718DE8F34201C1D018DD89616884291C14DCB0A3C985865DCEEEF58EB8593E1F7A7904E704653E74371F9C691BFA337A63C60CC1EC7F3FB0EB21BF8AD4E1029EFEFE5541A3447708D8268C70345620AFB46C5004D2C49996215EBC2D14302ECFEA6727A5D6BFD625FF858B8B0992F5B5DDADECD788777DCFFD17126BAF4109A74ED7A0E24E1F339DEF1E19C237D3CBBF070694E067C95FB08DF8C6F43B545DC4466C05E0B3748B3FF01742270F1CB619570E6EB8959E3E99D05A66BF2C37BEBE515AB6D3F495C397E636B9CBB9C111BF778508C73F190EA4CED77B8015E97F2F78EE087ED453ED48C6BE372452C22FADFA50A30BBF441FABF7D87698C6DE497F13723E3A5B6BE71783205AB2868CA3FA35AED4D3C73A0C34DD21972F693F0C47BA839F27FB406215DA997C65B4DDCE96C37EC416BCD378884831651D7CE60701B034C629D33C10B2F000134F1E84180AF6AD365B0AEC2D2E0A1B080DB26E9102CA17F82D7073523BA7CD0A8ADAA49ADD73F42A0B21CC6C70089AD15937F21B0935D77AF65BEA0CC5010874EB966BF29196100FFC274E359AD514ABF01B5FC21649B360BEF9B2A39034B9AE50DB4456B4C43DA6FDA72994A184D93C7134114BDA317B6AAC8F53D75D905F6EE49D6E7F5C48C6135B1BD9A88DA1FA35994EB775EAF760306B4915181BC51F61DF9361B6ED38FFFF4F0E66CB15EFDA30FF1DFA41AB8CC4515EBC7C2B47729261C1D08412D791354BB2431CC9296C2DDAF8982036E0B3A609651C53A2AA6E505CEA9AE27F02155EC21A0BF635BD63D9B145A655D48CF6E527698987FE67E76855D710DAA8BF19885DEE24448B8AEECF685FA241ECFCFEE3CF75E54E762085AC0228FBB8C87A2ACB57B3DFD585E8C8CDCD8EC03E34C290A521EBA4CE37B9E1F446B9F4A1B70666DC9705D6ADD69FC206B817BB73A87F4DAC204D1151E24B8FCF7F6EA0DD84D57B85FCFBDFAFF66C0CA32A0251D5CDF19252B2D685BBD746DD2A5E8263B5154838586B5CFD146587BB3CDD9F30F141B38575E95A7EC9EC0E4E6F412475863B9DCE3375B6677828690FB6699C1CC0C4D8290B5BCC0F500000000000000000000000000000000000A111A1F262E323A00";
    keygen_signing_kats[0].expected_PK = "D7B1AE0B7AC9DEBF3236824CA48B49A5FF417C11FE65C667716FBAA44D3DD620F5EBDF9D49AF3B711F815E9BB80488C8F3106EC723E7CEE24F1408D73787A54AD9185B8A7E331F6085371C71C5A94A64B11AB9C2C05D1AB0AB8E2F6DE7A10E3562C28D10C563C57517688ECFCD7D2C5103511CEEB38C17DB88D256DFB1282A2A8D668543C2A5D44E01419F2FE79A9CF7708EEBADAE74956B0715E9FEC122CD98163DE1B961A79C343655957EB046E13CDF26C3E24D625F751D28E8B08BAAAAA2FD10D8071CFE63C875E129B290B2FD263D306D502AEDF01423A182DC1608B392283D0C5A11EA510048EC026E3D53A8F6124BA59929C7DB8AD898A6277218738C1FA2E51B338E7F2B7BBC45F5AB90A911C62608B663FD5DBD157BDF4C62CDDC3A82D8C07D70C896B37B56CC307905BE965B17EE996A1420044941F3FFBDCC6398E3AC716C78DC558DB07EC6AB6B2BAE75F2C8EE5A27BA0109E1993017D98B42933D19D9E0DE56D743E6CC681E2179A6972DB9EDC51902E6527A3A9D7C53B66AF3BA37D62684C0CE046798EC4CCE74224A1161E8F61AD01D44814E34ED69A77413414CCD597588964CD1D9824E50BB818928CDCE1FA35D470101EFD1664AB86A4C1FFCB2E51CDF2072BD8BDFBA7440BD9CB8643D5D8B1833B1771FF48DC532BE02D57181CBF38BCAAC0302E0B499DB4176B967973201E21B6E0E4D5ACCB65F1DF56E3D855F7AD2DB23CD0F838DAC241455A085BFE125FFB2526C3A71DB0EA64E756E0A5BCEB7992B10518AD366DBA6031AE43F4AC033129BA2A206ED17FECCA6747E5F350E0791DD0656125E682CFF2C0176F6A6BADFDAAEA474702BB1A60B4169F506977C693CB34DBA3010A0D26A5E6C287907E5CA1714A93890D9913D86EBC5900682CFAA0CF01573369AF40708F3CC83DF996CA12530B54958A288F58CF0D95C61D5E689ED2208E4A1AE20828D1098F894578E2C6FD1841A583954B037B7DB54DAFB11E6D8F38A7A091D777B36A29F90744C11D4DE7DFDD37E9E494E73C2920DCA5D8A377DA84148F0836C88D472FFD371402DE5A990D3E374F9478B834FCA975D261E79F9024DCD70DBDA745C776678C17B62353CD93A6380B849BE5680B679ACB0113C004A616D8E3208F89A52264319F973BA345E16AA40825D14D30FB179E8EDAF525AF8BAF56FBD44C97E0A3191C4D9A3DB9D4F9291BEC065988D82D39A5284F435CC2BBFE76367AC78E9768A12AC88F268157ACEFCC0FEA6BEF6E520A3603AFC090DC7D922D779B805AA38FB31FD95D656EF5DF3620122CA83DF5E83051CBCC2E6767A9005DF0D65DCD0863A3B6DDAA9357BF31D9E370A027458E687F6FB159935101ED576CC1A1965B51F1B46856C070F3EECA68D55DE610111BD831D34CAB4BBA7CBEA57065E27C2E2A075D2F301BF6B795CDD8C91A8610DC72E495A90419E58BACDAB419DE6CA5A06498E6EA382EC2CC284DEBF0AC7D52417CA1310484EE64C0C8385839D66A48821BC099BE9C267E0BDEBAAEDF2FED4C8D5C8FA38ADBD77B153991516C444B5D9F7FB01EA442B3F603F7285896C612B9332DDBA545B8342D9E553E7AB2C88A320F9206F9C72FE3CBFA15EC12541EED585484D9E7E0A97B44BFBFB66C48518BC31543C680A7D320424BB0A22697FE255E4787498F998812C712CF20DBE71750472C51D4AC501ABDDE8B90CA21476383E861721554A9E667360E030B02563E51973AE326BD3F8B9BED05272845B9CAED94188989624D70FFE5C6758A6BF6E225C641A3B71AED6F2844778C4BA844940544D8C8AB1D6556737E995EC517F66A60B616BA243E1739CB63443011A91E704210637807B72A993EECCB0C9719CD2FD3480FE45A4B329E7FDF51CC8FE9D136381A2DA3691AAABC604AF98465EF36FAB8C2C71CB9BD1C6D48BFFB072206903C6A41516212ABDD40206583ED0F66AED210023B19DAD522ADFE6E31586188566B7C64FDA5BC850691C75112FD5392CB18E5B1C2A0BC79A5FA757C5463F134980F2A203A93F759F3FD3AC4A17C71C5C6E428AB13DA82F3A52F45FEF60C7277EE256424542309C371B33CA9D1865E9F52D839FA9E578187B6D0C7390DB1715596ED24250AEB7968BBC9C5B77A73BC9B2C777E49B73F918D13BACF546942FF5070B760C1E624DB603DE558787F6BDB326B3C93165AEBE0B818A943FEB8B2DD72D8180917B739789B533FE057D3154159B0ABD67B60FF681E011E152BE6749F296E778461277F5AFE8BDF28AC56DAC78745545E3C20C8639BB76AAA76500E799078E59650FC82A0CB2B28A05DBF574CD9A50AB041D494A389D4DD779814A2B24ADF580880E95BC21DCCA392CA6CF7E9A50A3D80B5E6855A0426182489090BB82F1EA2150016B4B3EDD9FA3A2F8D85AD61AC2807BD814E5462545B82388A2CD33F310E316D4815F8812AC924FABDABE7E696E0FAFF17546F359430461053031D31BF20FBEF05A6EDFE9720E9BF2DCFE15D83A597B3BDC52714778176C3823364B383B61F5ADEEB770C3D1FE161407D697B6201D5F5B1121D034A6157E46F81342ABEE5D7BBB8977F6209219BA4B8DE936EC87054132CAC3FC65666199F48C20E2FD56B08D04CCD4CFECECE2BD1C65ADC9D0B8F26E5DD582845B761350A3A8E6179105B7906EA2DF4CC3C21402F0FD5ED1854A11CB59262819DF514CEC51C026A2AB9481AB229FE42B3A0494FCEC6C2F6AC160742254DAE4E4CEB4BCBD288108A71805EE27B994BC919BBCBFAE1E3436EBD6AAC2A56ACC37DA6D39B52266FD3A6B1331BFE9BDEDE19B6227575662CBD6DDC5049E205F30272C151BC0CC00E3A2EC4A0E012FCDDE6C51FC33A18C297F86AE61803B21346040099BE7B5F1527E9D648426F1A06D8F8F74DB968D439C04660B8B14EA5BFF205E273283FB1B40B47012E718C50C7E899533E591B54F8D0631181962EF810298B0C29414882E51B073B19BF1C49A893E6B541D61AA48E2EC909102C954FF63E81C40B61BEA01D642B869002D6D8BB1DD28090DB3CBCF1AF7FD0A17108C3842C12B4B55B741C28E303863F74B6A1998D18A7952CA6F1A6F83751A5550EB32A0F9218ACF9945CCB1181AEC15D750B74E6A6B170A6DFBFC7A09EA13089B6906CDDD285835D841C2F27F380FDA69A0679FF94715861146C9EA97A728E1FC7A7AC23FFCF8150F94DBD64F47BE44207903C64F2645DC7D4963CA94D0B97E395341C8EE2D52D015446F972415A5B651289274F57D55705B8152ED2948F8BFC84D7DBB127F30ACF4AE91C05C8D5C964992A4E6E8DE6B569F4E36C5B846A85544916DBBDFF6C9250C91B9523D5EDAC17505D6BEBBBC8111E89AB795298CBA5A0E25450EB73DCDEB643C051133408DA8F3D6B47C1AE23F1B010473AD0A2F62E63D05800BF9FB05DDB1040268A0D4F0EEA7AD172EF547A9685C4BA4AC0D719E607E96D4D20314153A366029A81AB826BD5235228AA2230C6C0DE15232F7DF8330536A5A156801ACC2F20BAD0DA972A9FB2B4566B48F648A9F870DE8181484DFE57530A8EB0E5C214C418224699824CAE98FBAFFADC7C9DDAF635ACB7C92B2113480FC110E1D43B6DDE1A755C4E11F197E7C8CFA38195774B65DB88FE7EFE0839C22617E0FE33139EFCE9342D2CE72616CDD58D0316C1694";
    
    keygen_signing_kats[2].MSG = "9433ddf6e491cbf5cb03720b542e432f868bc7b5a0bbafd914f210c3a9d145953c6532b8212660ff219cb0bd283c6c25501aee58ef4201916e7671f92b759f21";
    keygen_signing_kats[2].SEED = "56594cac60a6f972e4317759f5dce7da43cbaa18717f89de21b83dcd3dcea9a5";
    keygen_signing_kats[2].expected_SIG = "9C5EFBD8FC4BC59259C5528538F9546FC47C6ADA017628AD039E841F3EEB41078CFEAFE6BCA288F8A1DBC40A0A8DD61D7CA0C5DCD435267B4352CA2E2F3BD346CC790FE55DF82A25C3F23D2D64B4A8970C1277A2522744027C90F0FA18BF22E49C1AE5E589129337505AB9ED4318F756911ECAB97C5E0343EAD34BA7B6B89DCC130903E9E0902941B58213C94C19CCB36033D514A628B3E99D819452A9298A76DF24407CCB332C55FAEC61CAB4C99D63586DEEF80323B8DC05EE160177046D298EBE7C7E07EE5570F6E4C95EA9F5FA6A72EE55FA7ADDBB09BFC096F6D544BEDD75DD1702203396E149C846D66B846CEA8A7718A627122ED3DA6E25A47887958A97A28F5A84A7B9E608A0D929CC0B48329ED824B2B39EAE56F20192F9BAC700C2DADB42BAD7210A76034CAB87576698AD61FC4FDE9A29193ECF2BD6FA5741143FF6D5DA8C125FA336BDB627C8ECFB327065C027408561685836107CFC2DD755E7933A2560B8CA5A13A5972C0F3CD1FABE9D1D31ED52E63EAB7C6F30D49911EE8435E1D58F42D24983484F62C6324CCA3AEF6279752CC429657C80E59D2CA789D82070CA167143B407290B373D5AE0F32715DA5040FDB844BB8B1B388E5131D5ED474004FCB10EEFA799CDD494397EB43DA9B69CE5468C13DB7E70E56A974B8EBB8636E62301161EE9CD92A61B9C00C389C784DC48EB29C3E3C03C13FDD841B6D5776583FFF2E143BA8279ACABD9B33B598CAED53EEF93333AD2076C5D4AC55625EE6888D67838B3FAE33068EE735F65BFFB8ED36A75071143D0DCDAECB0EA4BC1997778A6E919847B2127EFC49860DF42DB656681B115E7CA402D7395A3356957C9F63F6B53D7DD9AD681AFAD26A95B3844B042966B29961F2CAD3AE1B392C0F6E444F5F28F9D80302BE5AF3A450FF674ADEA63B72EA1D5E7C864BAAF1B1B2F6C65DC25073073AFBDE65BBD82C4EDFDA5FAB7C5639A5E79F4CA17143C4767A13AC4CD1942A1FDCE95F832577457FDEDA9FA8BD6CD91BEC05EA2AF3E77DDA26C233341147513E2E1E66079F6FBEDFB82B9C426516DE1AB27BC99C52EA86D16311AB303489693BAE687CA4FAF7FE5FF3E66D1B4509947C6A3AC8D2706C016BE4A75C64D0CB9F619B0E9310052D3A7DAA467698F54C043123316FB07CB095D389FAA0D643D9C68BEBDA18D3F26BDCF50C58271297F556C5F69E0F900C47E40BD22B9EC8F5762BDA9B6351817A93523B8C5AC863B8CA50E16798578F19DD85C80DD97ECF158944ED3874EAE1E4401B44FDB28053E4458B06B6A51C44635414CE5255C038FDD00B1777A12D52738298647E10B2C24A56932676305370B7FF2290D3907E1501CE17B67149CC83C19DC90BE28CD2BAFBB6FF08293FC2F0CA70B9083517F5BEA55BAC22BF1ABBB940E522916ADDACCF9B0BC1B2ADA06B3399F5908B6B517454FD84207A83C0813F1AC6802096DED339A162892FD2DA66B64C0E756360EA2A6D0DB794D5EBD44AE81263229F78F90543172758228F563CAE50C02B0E8918871D6F213A262B5C44D0EA31CABC478770B408A91FC7DB8E4A842E1C631951263BF836A338DA967582F4086D4A3BF47EDC57DBD6879D675322548705462912173BC8278FCAD7B546F9B9F73852724382A29F3904A06C8BC2E24BC0C6D3897A811A78EDEED0B8F8DEEE869542F936C7FF3AC0D67E55C95AB1C7A5F23AA1B989FCF97CCD2AE097A6E8548D97B0A76CBB2DFCCAB0C7D1AC9EBD3A8EB8F411A5712DCEFC79E9CFD3D69AF856E93925239FC666C7FF02518BABC50E8298766E953F95C2557637546DC7FA1B80E994F4EF93336122BBE707CEE4B7C2E875D2D1E14065A8636645A374D543E42586E4BBBA52D94E3EC1687C0488379A53C8DB5F409630586319033A06F7B21E382148906D16144FF8990B94FD90D4E85A729302410B89F121258033A7DA98883B50DB5E89CC9655CDFF8E9F041A075B7C742BEA13E36A83C5CDE0120BE9C59D50A0496A862432A82FC645D33C174DE11510873FE541DEA335E8054A0B193574CDE4E20CAB6E7731A1A28DED03844B3C76B9362565B332140F91AE84016758A0C4AA7ED931A509047A5F1F2E71DACC724808E8B30C96C5C1984FF406B3667937E7E9DA309B6A374DEE6E2C91CF7FD8F4459D4AE9D6C27310EDBB99390F897CC98D5A2051E848E8DD0BCCCC382FDB2DC8E4A4C1B5E6A582DA10C31B219E9670CFC53BB36EBCA29C6DF49E42B1AA34644FF5AA6C290EAC68938236913B8A8F970AF0A9A4FE56B2B441026ADAAA67E1BDB81D9FF9761D76E44CA7AC39B127048EBEDD8A2D41ACD9F559F2D0F575DBA0CAB52F8FE5E6031625DDEA9F363EE4CAEA36F4B6FB71CD079039867D22D089F4502A53B718A504F5CE1D0D16BDCA8860CD20D4F55A3D29EA7F7DB73AED014861A8C8E41EB39E3DAC98757EE6C3235673DEF318675D9E686FE85DEF0A3F38689751195460FF9BC8357191FB7CEB7A3F17C2FB1716301C5AA9550209CF8EFEF4A54E92FB41B1F962751EFE7A0C94B387F1DCD09DFFB76DCBE9B10D9436157C7B6755BD34321C99AB84335792EEC3730ACBD54E88AE9C0BF78072DF12ECD51175D4EC80EA45B2723BA6B9D4F5F7786A6F278078BC9D0FE09B4144FDFAEB86ED68A67609CE4CF3CE14B83D984007DA1986CB8488C0981C1D796B874DD70810601328E3CB1A72AFAC867022CDF07469CDFC1014899FE9BCE106FAFE9F909D4A25A886CF7EBCE107F52B2048A5D0A6ECA24532CBFAB0712B92EF7A2CB50EB15B2F9FD3FB0541A25E2DE4198202E9DB4B36012B2035F4F0FBC15CC6F121ACC19359A49381FDBCF74F46D80661996DBBE0D530B369BE69E0CA180D3CB9543AB8E7BA2C7BAB67C7B02DDA2BC9D070A60655A9FB0F90E6468F7502EFE170871FC0E27D43C3945A292BCF9BC01A3FDDEFD87E4BA46D915D918622998EAF3F64C3434E39B201921811D67F99F964DA3A831D6407F1C8C5311557E6D9FB83D55A03F19E6ADB056A1E965D90D1AD03F9B8588DBDD78FCEF81DC190944AD7FF4B9D1ADCBA06666649E5D8276D513FB7E148F3EBD555E0361A9D204202BE359BF4E5FB7A088C472EB0268323CADC8D5CF4E74BD9DADEF65A0395C26D57CCAD179257BBAA1C4D39B755CD3552C2A5A0C53ABC114AF180781F11AC83E7A5FCF7FD5A977A6223F6D779D2982B1E82CD6936CE4E29A6C5BF88D474F6FB163C6BF54F8C19FD556E368E71776048FDB3BF51E54FA2814DEDDA42FFC48A00516CF304CD8C6171922BAECDCC8779B43B73D8BA39E3C04C22745C61B7D92EEB8BF28C202375BF9B8801408F036685D0F04A11E50969BD235412443C4503560922750CB2BE179E4C9BDA51FC290ECBB5F51BA7CD060F6EDD70CCAC48AAE5E05E070A01874605CFAA6A5844B3C20AB989F6AA03DC0E9C5D046EBE0A819DD770849BB0039A1600AB455F46A0A6E11FBFF35CC06B4A87099B07F7C62997F0FC4BBD46F9A0001F031B58D2C1AC8C1B91ACD3BA2E3970B1AF0D11DB275C898A7A340BF0820F81370E957590F0E513A0D128325BE86C84BC61815BA37136BAEE6F94E0D0350758DF89B25CEC22D36515723C90B697333359AC830D4CA418859A42255163761642B84704DFA6E0C835560BDCE67E1D5424876053BF05B7B8310E0BB46299F3CCD677F8C67596FA268368463870DDD7F06347E8BB28BC7E3EA10ED6BF20A6939225DAEA03BF52D957990EB0A8DFCF403E67D1EA6EE6C48CAD03580883D0086546A8ABA936BD6C837E07EBD971245FAD5213EB5CC73AC6632051F5CBD5FC35F143BD8A30E4CCE9CCD9514626B986F2AA0787CDB0CF797623C41C6786A4D8F39C6749EFC1F06E968692C8B67ED4032200DA35A1C2CF393CF1851A184891F15EBA55560D12EDE777CBF5F95AAA638BE56977A0611E004C82ADB6F95906A3949BDC01683988348D3F5A47BC0BBCE22F7F147C429EB8B9E2FEB013AB6D20562B3E2856D4767AF8F8DEA16FC75815D9D25AC13795BF976E41FF3EC1599F36BD913E7E2D9AB5ABE7FB6FCF2CBA652CA00C3D84DB05C4BCCE42735822825E3DB5580075CEDA00F0F06500413EE11733C8C1B7B14680FA368EED79F118BE06E8373168B83821A2EE66349473CB0C36B16C4A00EBF9247B9E187E8CB4CC2429F3509D91875CEF69AA95552299EC7EB7947D6F1AA41A87B8DFD40F4F3D2465D7D1B26F0C4568448897115C4C3D007EB35270AA60CF47740F193A920291ED247FE5C67780F510FDC23A16DB4D1F56E4DA799EF2245BC2EBACC2D6B5564758F33A81E1BEB3075235AA6B132BDB0EECC4F98604138700D3D36C5B952F84CB50820805E8DD2D46E7ECE54B2EEE4025E158743C0D9422715ABDB76934237BD743ADA2795F5881B1A4139A371156C05830BB656A0D5571B419894D52CAD68E03C64CC33EE70F90819CE89A91CCA0F5ACF1594659DD195C8140E02D0249EE10BAF3C8068B765188627DAC302ABFC5A0B30AAD53F476C8E8A201CB5FBF85055D727894EFB3EF70C991A2D9D6C411923E456F4F8417705F042E890AD69AEFBE5E9EF5C0307FB1A99CE9E99C7830A383AD703503D5D847D703150920C423BC0A2CAE2A8E16F1FF30C932240F5B9239A4A3D4E56AFCCDC3A06E74FD5930B336052F9BB6029AAF9C9718AC62FF8352088CC6833D5F97352B4176463D58CE514D458CC5EE2B99E84CDB24F760EF7C737FA0F762FF4544BFAC078D4494C0BE2769EBB872802590E21E94599257E9452161968B6C2F8FCCB8241A861CBED00D2C38C3438A8A5BBC44C533B9B8BBF6E4F9DF7180BEF52062A465BA266B97021D16BF0FF8E29044F1D13798F47FA12791232E969484F729C699F7DDEFBE97E5ACA8FB900943E2EF04CEF3923DB07B9AD1D2880656BFBB365CFF326834F651A9A72181AE1AF6D9DC7FDBDE84F7D271984F948B8B963567F548E6E00C1648EFA7514E072C603450FACDA79B6827ECCDF9E607E9B2229F4976D5E7A3F3E1415854F2BE29A585B23FEAB97EF227BADC65206F8325FCC362A00AAD7B8187B61BE1AD29970EED3D6434D34AA81D6AFD4AAEA7CC5E74B43433FACE7E078ED44F84008D7CA3BFC44DCFD87E27F728FC2C7CCED887DC03D875305E266FFD83CDC31FBD75D17D94192BF7CE72259C37F83B2F47AD244A77E26B07B014A5F45003A433E1703E850D6BF96129079BDC684EB34081E43BB2020A52FBCEC34C9F035DCA3A66B152849D34B8E5BD492E06FB3F96145C52C56413F68101E609C93DD58362D24F4C849DB5209487FB47CC05A104C6E55E4F275A66ADFF772C84BD9B5651789982205367085DF95EE12B8CCC0CC6E442F98215A5C37952A732DA0E779333E1D35F75DA0F56162400BE8ECDC67F554AFF2A791C7B67859F1BC913F934A62CBFEC106841AAE74E88737E9C2C26305A32F5D7289BF25787C3C43909C175F40B895F3D8E34BACAC56F6406AF5F3F1AC28707099F68D72C841417AFE98F6450A46FDF89DA5909A3F1AD6CD16D6530396D991B6502D137A13BD91ED9A9461BDAA264746619FB4FA93B843580C68AAF80AED82577D16CC4E354F9D90EFE35F0A45ACA7D39831443448091B7308164D49255BC12FAA901E7BB0B98664C58B5DEE3820BC3497F0086B8346885403502886329442C71E51F7BC2759DB3E93F2193F74B5D923C5278D1CB41B6943E7F09FC36937A7E9DFEE6D5F20AA67C416123B66E7BA8E370DBC11755F912B65D16E29E4F3EC01ABAB2CC40BEF9286C7565806815824C3A4BA8BB3430D4DAE5EA46EEFFDE0BEC592EB00776E06D29D76A7A8ED633429574C9F9515C149181B9BE8489840B486C29213964FD8058497424832A4D221964C344AD9731849B654D395C18F2117CC3DF86B8BB37CA65BE7504A3FC27C9EA0EA49893BEA01028751C51826163AA95224ED6FD7152FB0ACB25C38017EA5FB6267CEF654BDABC122319D439B6173DE4538DC5118269CFFDD446351E74811FDEB87D3632C4D2EEF56AC06AD5B6C339F15BCC6898E36DDAF4B6A5ED83C37ED5C0B9E67372C1422302F9089452EEF0AE1D53A81200A44C6856ACADB838015B18932E682A6F7B2FA6CC9943F63469AFC460DAF780A472F31ED748AEB194CDEC5768B1B343AE64AD65985F84B5FDB0C98BB231B86D99DDD9C1668AE4F333450A713AA35FD96614EBA5EB3400681653327698445866C05347C84AC8A265930D486F08727633CE13FA0C844D3821F5727FBB3200AFCD51302E199B80F4447868E425961B19C8D649057B4FEFCF10EFB016670503848A1909868460E6429C6DC725E2FB5A73006F929D8F71DEA23B527AAAD638180E4339E82C9AADA5D06B8ADD5BFB077184FA270854B613A639084E6CBFC6253011D07F8F045CC391DB45CAE21DA014B3D67B9F55E6B04212243577086949CB71C1D7A818B8DBCE818254E7E85899BB1133235518B97D4DFEBEC036BACCDE0F6FD010F687F929EBBCCD7DBDFEB03579397A0C3C4D1E60B103D8EB7EA00000000000A121A242B37404600";
    keygen_signing_kats[2].expected_PK = "58E3563D36F5D0492030B6E5AA317FD727165ED2F494FF5EE45F7E395045C87E4B5709DFA6E7688B11B81F70BA940DFE52729C62AC9C8D56B0A93D2D2EBF4347144EFBFCAE4BF801CFB1BB6570A8A58C27602F44DE8399E1EF6281B84DB2614F4DE383BCF4573F411FF97CA729BD3503FB2F91F5F778581E89A8A44E3C3C3A86893E78F991B7A7FDADBA06C938A8FFB66F58CE9B584FC5DA89190BA94E896784834914A4240BD8143E1A12BB78036168B09D1E4BD274FEB8084EAF2913617D2A1C6BE16B54224C552B7D410A831941EB25AB9ADEF774A1F73FCF1436D428E051C23B2C7B08CA788B5A70768FE2B6B202139177A153867A236A9FC9CEA37F47FB7E2FF30972DE89C0850DD7B38AC0F855BBE607FDCEC0E4A32E7928450EB1A571357AB0E137830379F9BC7AB2D8D25C3C59E56229A4DFB1B28BD9B7D8A0B5FFECFBADF3D24EE4E15CBF34D6E771AEE04CB3EF866083FAE94A7BA0853AF896B1438FFA79079DBA05ED1326479B79EF1B770057907CE068B3A62170936F42DEA21E596710A0975BEBB86D605A8A1A4612E47F9E60678602080C57D07451D6F207DAC1D55444892DFC4783FD0ED05DC61054D1E5E234D11AE559C35EAA3A5F6F2EAC9F908600FF2229F188B3C7C3488C88C891A0016198F6DDC951DEC5BA79D217A7779D18938536B8A049A8E418E1A73B77490A8A11A7FC28F100D3F706EB490AC59E38D39F30BF632B458F4CEF494D5132D6C74864737D05AB0AC85C34C91A19E4BC065EFE5BB4F27718D9FFA0431E5619F447CB8C92111EA5AD8104C57C47E5BA02985D0DFDEB9BC9A6FACAAF57F4BE0BA680BF83308306BA43838F7EB9A8ED5F1384134902DE002705100E6785B2DA943ED591CAD0A085A850838E10AE9889FFC1CD2941E1899E1A26CA56CB7480D260B217798056D35EA62BD55F159CF0FC363A4F325235ACC231BCAE18E89EB70A6970B2EC08DB004961FE951F8ED294D7D68CA6DB402325D054A47D17FF5B38734298B99278273021F165817E7805D581A0B9E40D507CC89D543F7A1B718820B1F8414AD6946B1AF7BC3AC1A520312240C0B499CF6B2742508356F9C366980BB1894D343E1BB24F06EB81CCCF5CAD59158FFD2C0D5E0019A839EF8AAF32292C33E32F6454BC03F7CE05D157BD875210A4276EE7C828291BD5AD5D545AE4711FF0C1332AFC7D716D104344E88BE87124ABD94216405A370AD8097D80879DDE60CB1F70B8F2230CD81D719EBF1C5C1D6EE965A85CB8C9982CF1625BC69B0C89D5D4207AD037DB73A929F024DDCC2306CAFBA0FF819CA596EA988A366901172C153D7D2A467FA1AC7E738F3335C1A2008181A8EF3064227FE7E72DACF26BB28816BBECFB8224167224BD37C5B55BCBA256C9CBE8B18FF4C36EE6A1EF091A714416E91DB1D638592D0FAD1DA51085D36D12B1255884B849B2B6C661A9FACBBBD67EEE7BF27CEF998FEC1CBA2E5EBD5361B429D509EBFC6CB2DDEC67B6DC69884A342D4A6C6D8001E9652A1486B5360A17BBF3A47DE94D1A32A5E2602FAF1A41B5908F67E9832382E87C9D432A3B8B6E230A58EA733F980488491E7043F327160FCB6D34383FEE41FE7DB76D5BA72B3DF23034E648E8ADAF8D53E1F63403A62CAF6AB88CDBDDEC39E9AA4233E3D335DC890DB9454CDFDED997B292562B5B001451729C833627E9FAC08097FDBB64464CE6B4C0D33FE64987373951F2E3E19E7CE119A82C2529C244BA56C7BA3C703CD7C940759403829A505A635B4401AAC9A8A9C76EB375F6069D6C3FB6511E20F1E9F1B40EC3CD47CB90B638329F17E1A3D9CC45769AE2E6CFD9284C11F4B0892BEA676F9B09CAA8E83CE7B7648546FBA7E7A8B9580ECCEA43FE330A0F1520F5933164F524CA22EBA3889A51D184885E515CEF8B35E65DB4DFD90D8D4FA1FBD0F7F0936E55643905AC144175A27F189865C011D8570E2A57392A521C6C38DD7CE0D3FB5FB4C34FDA41645E5BB32DF8100507B8C0B33846D12C5878D5AA05B86E4D83718B5158E67B4D8CEAFEAAD3760599C63A0594B64E21DE4C1734AFC875005B798550F02D1203D94202AF189F140D3729733C276DBD47DBCC0B427CC113A38382E4044B74333D6EFE559FA327F9EB5DA8CFAA99B882EE97280E7A909E4B23A0D35CA8164440B71699D82623BD542ACF364C6D74E4D8D79A0C293629474B5D8A05D3408423A17B9045E9A3A6245D4F123DA541FB8FC8C5BFDC3E6BC508B823DB3EA81D1529558416E720346DEC470E5A7FDF7720893EC139DF5B8A7664ABA3FDE76AEEC0EED445850B5FE0F81FB3D0CB9BFC1432EF66FB8960E4601B50FCF176AAB7AE4C0E9328CBD5ADB4D8DD89DB72B0221382D96C04A8F511659D62FB268D781EB68962D2167806C73916CD66DF16E9CB7A1C25C794953FC3C87326AC3195E6285FE5076C35A56F24E7583E985D51F8EE8CF24AB0E78F2873E426C20B94D15A1E178F22D96C4EC22E90EB07EC066CE4A19BDCD66D03CAC9DD906D9D85C630A7E10F118D83DC7618AFECF90F3CD32D265253A05FEACD7DA610FC868BCF54F0053BB7625CE2E2C35C8A24BC8F3DC294F60DF8F345ACF03B2D8BE69B36E51B49492E8891FC09787527B3BEB02E6B2B69158448AE4507FBED5C3FEB923854656B642CBE0176DEE52B92EAF411B5E1480738476037D52D7AC9C04D909EB7AF11D98BFC66DFFE81F19CE1AAF2E3C646679B834CE0030A6E3AC7BE93027D2D7347B9165F9DEB26CD54F33A90A3AD5FFC88044202208C3D1C97B9668542D6F1DC4E1FD2DB6489392E9ED43FA989E5CCD6CC63E357D516167691AF5558541513B38D8DA32D19133EDF12E1D161C5873BB423B4E52D6B34E97875186D0DF7BB4EF4D05023B19274FB1DF47631F6282A45FDA95A07F8D5B0B0F814AE31CF30947FFA65D940C88CC191B3DD031897F8647D0F8D68C2FB79050F90EDA905673B206E6BDC844875101AED46513041695E9EF151B06AF764BBCCA82B0C93B9D26AB96877B49C9368C972E5D42E2CD41B3F7AB17F8F0B3EB1D0C284C699D9F5523D6C5E2F1E33747E49EB675CCF1B68D2CCDF4C7CAFBD6B1254C141001BDA1E8A9FF6F05C8B914182BC4348655D69D7DE203ABB70242AD8851369AF610CAC22E62A9B300F53ED948BF17D811B6C6B65F2E858E645F95A7F2DD7A9A6D6C2D627BDDA4C852C2AF523F9D03109335639009697FF25A1C67E3100083BD6A741A5B4C8D5567A85820E3D9CC6A7F03A1B7C902C75EF1DC49566A0E3A12671097F086CA024E61DE92F15303B0D6613EDF5FF80A5AF17FE2613437263899D8F66DD19B34A7887B72F416B8DFF7498EE37590DE4B1AA099E9AFE8B78D139238AB3473B60BCC70616F6ADEA0CE912C640D4672C4D68F2DB405ADB6643D7C82EF4F4C95DCE932DC8C96C870B1B7C0B91CF5150EEEBE6973068A3E60C5DE142C96A2DF5495E1CC3B3823608116D0838A5DA3A8AEB40887C08E58A62EA753FA3DDD0BB615646CC2A5B185C7B55A7DDFA9704C4FA0A74A2B1BD579C24AD9110B103A6042DC329CBFC728152533A41C3DD19C7F07F5DE5C863C97DA162E01FAB8E70DC91996897C68A173610B61558F298EF0A540BD762754DABD89B89334A2F95A9861879E0D23DFCA4DB8F04DB6A7E6A3D67";

    // Iterate through KATs and validate
    foreach (keygen_signing_kats[i]) begin
      parse_hex_to_array(keygen_signing_kats[i].MSG, kat_MSG);
      parse_hex_to_array(keygen_signing_kats[i].SEED, kat_SEED);
      parse_hex_to_array(keygen_signing_kats[i].expected_SIG, SIG);
      parse_hex_to_array(keygen_signing_kats[i].expected_PK, PK);

      `uvm_info("KAT", $sformatf("Running keygen and signing KAT %0d", i), UVM_LOW);

      // Write SEED to MLDSA_SEED registers
      foreach (reg_model.MLDSA_SEED[j]) begin
        reg_model.MLDSA_SEED[j].write(status, kat_SEED[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLDSA_SEED[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLDSA_SEED[%0d]: %h", j, kat_SEED[j]), UVM_LOW);
        end
      end

      // Write MSG to MLDSA_MSG registers
      foreach (reg_model.MLDSA_MSG[j]) begin
        reg_model.MLDSA_MSG[j].write(status, kat_MSG[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLDSA_MSG[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLDSA_MSG[%0d]: %h", j, kat_MSG[j]), UVM_LOW);
        end
      end
      
      // Writing MLDSA_SIGN_RND register
      foreach (reg_model.MLDSA_SIGN_RND[i]) begin
        data = 'h0000_0000; // example data
        reg_model.MLDSA_SIGN_RND[i].write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_SIGN_RND[%0d]", i));
        end else begin
          `uvm_info("REG_WRITE", $sformatf("MLDSA_SIGN_RND[%0d] written with %0h", i, data), UVM_LOW);
        end
      end

      
      data = 'h0000_0004; // Perform signing operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h", data), UVM_LOW);
      end

      valid = 0;
      while(!valid) begin
        reg_model.MLDSA_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLDSA_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLDSA_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end

      // Read and validate SIG
      for (int j = 0; j < reg_model.MLDSA_SIGNATURE.m_mem.get_size(); j++) begin
        reg_model.MLDSA_SIGNATURE.m_mem.read(status, j, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", $sformatf("Failed to read MLDSA_SIGNATURE[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("Successfully read MLDSA_SIGNATURE[%0d]: %h", j, data), UVM_LOW);
        end

        if (data !== SIG[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("SIG mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, SIG[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("SIG match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end



      // Read and validate PK
      for (int j = 0; j < reg_model.MLDSA_PUBKEY.m_mem.get_size(); j++) begin
        reg_model.MLDSA_PUBKEY.m_mem.read(status, j, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", $sformatf("Failed to read MLDSA_PUBKEY[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("Successfully read MLDSA_PUBKEY[%0d]: %h", j, data), UVM_LOW);
        end

        if (data !== PK[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("PK mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, PK[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("PK match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end
      
      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end


    `uvm_info("KAT", $sformatf("signing KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



