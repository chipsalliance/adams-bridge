//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//


class ML_DSA_verif_KATs_sequence extends mldsa_bench_sequence_base;

  typedef struct {
    string MSG;         // Input MSG
    string SIG;         // Input SIG
    string PK;         // Input PK
    string expected_RES;  // Expected Signature
  } verif_kat_t;
  
  `uvm_object_utils(ML_DSA_verif_KATs_sequence);

    
    // KAT arrays
  verif_kat_t verif_kats[];
  bit [31:0] kat_MSG [];
  bit [31:0] kat_SIG [];
  bit [31:0] kat_PK [];
  bit [31:0] VERIFY_RES [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    verif_kats = new[3];
    kat_MSG = new[16];
    kat_SIG = new[1157];
    kat_PK = new[648];
    VERIFY_RES = new[16];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // signing KATs
    verif_kats[0].MSG = "fc2925c28f99410b1f0185546e7219797299369d27c6ab2d00adc627ba5564816fd47ef3175a769ae51fd160d23e458403e27cd6d16678ca6367a098d62e6610";
    verif_kats[0].SIG = "277F05029232D41F8597688093A174585192D0CFBF99ADC0B2F2B2EFC34E61114B7C427A0E05C24FD7143FE66213225CD2F0D707B3D40F17BDBE0CA72D1EA0AAE75EA1DA1E554829342D1D83953607150C60B7635282298AF8E46C0E72CAB64C52BDD8FEA8AA243EE25531E31FCFBA93BB298094D472261769FC3FD0DDA710B79588947782B8C0873F26753373030FE87A6CF390E81E16EA194162F94D645CD2A100321BFC008B0C1CC17C119E3F585BBE9187A5CCCC73659852D236E9A6A1886012986AD3F3DFBEB7DA0D7841CAE598271924306DA59647B1083523CA536F4BFAA2D8C73FA03DB53BE2AC24644185CD27D0904EF1F1DB2356062F93175D423ACDCEF9095E46FE14EC15D128A974C9551F5F84CC5DAACBBE0EBAE4BF5E1E2AD84173BC0AE4869F9D019CB35E6483BB3AB793CDB1C38287AB1A231D333A09E7BD546D696485753F9662EC889B62FD872926F7D79FBECCF400729DEC7478BF4348D8D572A2C78BDBEDE62F93FCE3FAD2FE3EBBFE55EBDD57AF8F2128775CE37172C08E3B3249818CEBCA291FC81756ABF06853AA2628522DD1AC2BBAD976E37C30299918C24A3DC3C9E36DA0D8FE6CAC8427739D78541C89A098809B6C03C002065B6516E0BF06155963A3E7EEB6168293745647CEC9327A2466E56018EA0C62A2F9C40DE2296FEC58EFC8D863EFF088137E0BC9BAF3F931AD163A01B1C65512EB8C2CEA1A98261BFDCEB9A28A77EF25035EF99569D9A830C51F7428545BAB1EAA495E788B3AEAEE7EA0F7245CB3459F9D57711B15F8081BFAF05A991A3696AD1688A108F38A16402F1CDDA25075A2F5AF526DE382FA337288BD08480B46C80B89D5DD93B2FA5AFC6D98016D1CC1BFD91724689F5B648D2748AF0817CA39F176D8390D3BFD61D1CC9D93E280E141C7F4D56BDED7068AE80DF60F19B13DD916B5BC0D7FA974B27D36DBFEA2CABE557C72CA39369B216067053E560586E27E93E9D15D61749C6A55CAF471B7DE782893642D7B2AEB83E319F159188EC232F32C14F5C43FE4DD860DD07BC655F21249549746B6831D75EEAC2DBFA3A9A37752E984200122A38C1B3259CB01BC4A3D9376EE8B0DA134CDC0D475E8AC4DA6D38FD1090C2CB7E9E28AAA4DA7A396EBFB1E268A6A1F4224D8E30F9F0E99468E6B3E416CF1472300A245EF25BA7430B0039A342D8B13BFE22296A01A3CFBE3009C652581BEFEF0BBE6D72FF6479601440C91DC4038E30324D942F51DB5D6112691BF00338F8EA3108AF6BCADA13D3AA1D65589658E51432C22442B02E2019696DF0472D6413D895AE3AB88434F1C81C45DC2C0858D5F1843E23F465C27C237F6F44DB2BE13AC7C71F9761AD6700F9271A3B9CB93A6D7D17548FD9A0C7D696308B4D54B9761FC96294536D2310F3565764A4D0C8E3ED79E9D1A270F08363D3169374645F63C0982D4324AF7B2B95FC08A76F93F66FF675C1330A27BD577198D2BCB23BCA01FCF62E2C6028CFCF18CBA98C3F9673A69F09EEDA06BBF3A97EED9796A3B58F279D0331D751F40755058F6721E14C354B3305BD90216DB2B8B9D9499DE8C159D4F9D22925B44D2B31F291C9EEB29BC2AD5E8CD4AEFFC86018DE0060A027363E67791ED08A8636564974BFFD02CCEB42C91788374CB5660AB4787AAEDC3395D50CA94A1AB7342C390210B48CA3EB785D63318E7F4224ADEC3D1421A388BC1B60EC089073F40292009CE51A010F27AB94FDE6EA497FC28276F3F2C3F1E3E22177F262A6CF581972DD5D49D8DE3A8B48D16B393F6981D62CD42AD28166BE10FEF43AF5D44FF15F152FDA66F46DB34A3C202D4147DF514B38F3979682AAE97DD66C4D5BA343F02B113508B4668A64D2FB549D46533A4353C5927BF6B193DDA90EE6337E63C144913C0DD2ABE70972B2A5160FFAE8C51767F0F77D786364F60AF4108FFE5848A6B7B7EE0DDB5810FFDD6FDE9A478E0CC8003049ADB59362CFB05F9D767D3922E620BFCE53BFAE26FE813B8A340C59125B579663A07F1015E9DEB7A0921D79A9A3E9EB4975C1913E22F0574CE49DBD56178157F46E3941047116868A2C79D85BB6FAA3B55562DE86E12EA3AF24C4746D79CE96CCAB8FB087F16AAD2B12058721CD1BDDF52E3C1EE0A1FE129EE3D0E0485D9D0A1C7E2A939DEA764D88E71CF0571390F99FABBC495C09ECC3B0F0B09A76FE9129078A54AFC5DA3CE3382469BB962731A96A38048FD0BCD70BA077CB3F098999535F0DBD8F610DDE6CC21DC8A0351DBEC04A3A16C1BDBB70822F18FB02A356A18E496F8C4F0BBF71330634248A04E947C6761932F0250C3DD170E976D3D60DED07D78119A106793A1112EC1EA1353AD65682A40C01836B1895798716C7169C8DADB01D11A18F15DB967185D45D5B578A1DDBF8DEBE52ED5D6D8ACFC555A8561C6B0D86A4924CF15609359642E321D59BF8B16C5A22930BE7E16173119A2263F48919CB92A8173CC9DC10734B95A73E5687FC27A76015A0F5F059CAAAA0AC31FD3864FC26D09D7B11033C72DE5D85282BE3726DFAA8A1461B008A7EEC42081E0369866DCDC68754A18A94C5DCA1C635F220B953170140B8BD7D1705C951D0CC0C42D09BF7B69A74602EF55CA68B4D9E33B4D4C659F2C7342896D7E2F181FED0868AF4F1BCFF04C8E38D7658A7E000254C41BB4FE9539DFB912DCAE5807A35677AA72EA74E68A02D53BF786AE5B4F09C115058499A7B17342941360A98DE3CCF8B7E5B4DAA70E80A98A34B8921E396BF3F72FFC67132ADDE43E564B3532D5F29A65292A558928F248FDB14CD9FA553E81EE88776B60325DA56A8EB800C5ACE397EDC1C7E46F2E2038527016E72051DCE217F0B8354F9B36E18B5C687997ECEC710406AD27D7C9651871211C76CFCB8DD761844596B873BFD3E58882A72607E36173318D79DD6816D5CDB4CE5C265B86A99BD745BC86F121FEC06B02D14ADE60D1C56E0F2AA2B970D28233124071BF25D17B6EA917B7F52BF19CD6916CB4AB142C90C247E8FA23CA766BECC02A3BAC77A0935BA8F687B8EF4A1895FEBD68252AA32FEF8B9C9AC928C79C7ED70BE4B0071115718EF62CE2448D34FD13D57E84B44D5F172830866C7939F0049F09A1CEA9D908016BEBC54E34E08E7B7D8DC13E45456443B29A3694EFB0BC6F91242D38A641D6B49191A87A2909BB9339AD0506829CBDA2A8288AC28D6830DFACBCE5BC73CDBFC7B80C070F1C3763FA1CFD03C97ADF2F3D8E1E3A48223001590BA8EBF6D9A41B2B97CAA9C8563B89062B9EC72A5368A31F25A7F84AACA334CD932CAB8CAD1B7D19F5B11141EA720DD59BD719319CAB3783B6C0A99A0B6CFDCFD9E94FB8FB9ECF7DE7D5A574874AE8CB1D9D85EB52B07D886BAD908A4CE4B23CC7867CFDAE80BCD5FDCAB03D0BCC5911C717B0C3DE80A1D1F97AD7CFA0D48C217BA6145CD26925D0E82077438BA442AFB0A0F246657724D493C3454A389C18626DE2DEEBA87968209DAACCD04AF249F8EEA09F85F3AD3CE2891D1BCF087A983E20327B83E60BA7A0A7304C9B1734959E6260D8725EB71BC039D9FB1B3A59DD2C92C9BDF82AA091F929CBF898F02FDE1E7D0EAA65422821FA516E01E9B6F9A23C5C4D9B0FD316E2D221482DCD2E3FD1AD8501E23E276CBF134F039849E726C51C1C4B3D8252E48AC4FE2FFDDB5EDBA472CBB4DBA98D5FA859F5DB814E323CDAD0087454E15CB057AD97CAEC1BB346B9D77B7C35D1CEA1A1C1C950DB2C29807EAE7E693C844CB3731AC26080AC47D0192C382B7362A62F89A4D03F787BEAB7F6F60C4FBBFDF771C69B8632B5DB955AD1955C6C5971C7C8E38559F1C23B2CD95FDD53F4DEC0128AFC291B0C15B845B7788AA645ED6B27BBAA39C052A611AA922D748238583FB8DF9932ADCC325EE4C52C85D24260F680E71F885C70A136C6B7A0375D7FAF826E37ACDD6B60915F294876E0106E77FDA6DB08516FE156A370C005E492CA5164C6F879D2E5ED5739CE5F78431FEE2AA1A2F07812CB341CC55A3D963DA4A64821583A3EBDC0DDF08170F98390B55D571D474C9C68DB5F18FE6A593D6149351A9EE59C21E3C3CF2E505A07F14202CED73B589BBD44626116743BF8588A9F015F6467F09F511AE67AACB70027F7308058C4DFBC53775A78C80FB10B723554313C3CAA9CD8DA378EFDBDECBDB5B4F217AF6495622B85404A9E890F4018B49BE1DB706A4F3D988749D193BD650CD6F83761D269D1BE13D414DB9C7B6AC6893822E7ECE6B0B05F7DB323F65CD51619BE54E61FDF727F885FE8EB3184A894C7B907DBEB89777B2E744779729F0CC7249FD062AFFAE7F2844A99187C7233C71DC12DF657C92BE221489CE1CB86B1A1DD28A549D1D68EC33E2B45451562A278C648F94E3E971BD63CFB02D875EB5FB6BA8E4B83C9EF92377237F9B16D0BF286A37F561FD53C2EB7B0E6D12468070F67E69D1C6D96CEEF791B3072C083D735BBDA4D502B584234B8393F14135C688297E54EB05B811E9851C7B47ECAC8EC8D9148E3CC0F365F2D39A9F4D5C2463DB4C7B5DA73E911EB643FE99A517F6B0B0803EA4F46E663BD1A93C5A6F3D1213869CE001EC0841A2325CED0049D601F9502A74B290D3952ECCBF7FC0981C0F68FCD56BD7964B9CD87DD1B3F6D5D12AC536741112C58548BB110B15339302B5FD5D6FD9D58186BF8B788BABD28D67D5E400FDE163736A999ECD9A112B4BBCC320A3B11532E2D24C2C6405651C1615B86009911F1974E1A53C1AA7F0107795C910D3986B6119A661A19D3B62D3CCF415046C43FFB9C72CBA29DD3F4120F7B8C305363D15F0450E5C2FCBBF5AB8CCEB467DFC426220107C452A8A5A3B5263C6138C1C1E910E064E8AC2337CFBD9C11E82181867F5733E2433426466D7E7E60FE63B6C70DA6BFB515DDC0295E807BB6D54DCD7402025743B2F9BF53336DC3B5CFC48FB4DABD8CAE2DBC8043D7E57D90ADD5344B9392BAAEA0C490840DF046F0E543BB56F33A7ED39C0156077174916F276CC91007861E3675F4DB91B05B6AD49CB5D49D76FF543FAD37ECC70E81D2B868A75FB3D72DCDC3CB84E993715C987E8D4E35AC170B94CC30BFF511DB46250FAA39FC721E6A877D5459A91EA5CB0D9AD3FE5ACD4D99F47D48CA718B2E84A2CCDC187AF464052D0CED4D665F39106519D7DF9B345C3B96B9F1641CFCAE0D9E301BAC5BBD70973930BC1FE6FF9C0A5A5BD4C1CC0AF6377E3C6C267DE6EB8617537B45CB150AB5690CAEA3FA2D3B52A7AC4395B39FCFA831CA29E718DEF50D8620F97E8B3E95250CA4BE8F0B9373814E837B43AE31F55057B6E52B8775CD42E8E0A1FEF90A25C46A579D9129797D8D0B291A244B1EF8CDC4CE6FAAF327587C37B97BF2B6B876A82B2EC5E17C526B8306B632A515EA475D351B36D088CF390EB89CC3643008E9EB6599F845F82CA7FD667EEA98695A51AFA7D1F7FD2463F0EBFC4499DB3FB07605C3F502C42433970DDBCA1791DD9920AC9876401D30952C90AD1CB3542E13FFE0F88170964C8C56ED03CE9F2F40C7AC546794F5D39263D9C3EEAD8F872E830225CB28170CBBB6464F515E7EE8090791CE944521155374EE6E544E7CF5C15D5CF61F691F6AFE6CDC3F243B270337D436DA06259BD3091D7D4298F22A126CF5B0EF27D09AC3BC8D472E9EB6EEB1356E69CE1E7041E21DD09925E4C0735D7E00370A09CDE04D93B13707B7C52FCA7BEC9E10F53B29E56721CA9CD80B28CFE090DD0E850B11734691B78C335F0A236C9A3C7FD349F6943649A2DEEBA09EB0E2BCE86C76380440ECF67EF30B622D9F96696E656ABA4051727D741189BA271E04FDA9158E60E8F93AA0FDA6BB590031673B22F96C2E4CEADF52903FEA84806659C7E5301952A88A4964D0BE4BAE39251C2CEDADBB70D6820B0DCCB10C20B570B20CB65E25441A85C99540656DACB6580CAB798CE64A5E7A2605EB36E98B06DB85B486BB9DD840C05D9A74805857BF229DCE796242F8AF2297305E595E933C7183D475E99E38A983B5D779CA2B6C2B8D1DAE7327F834ED2D4C140F94DD1810783DC308333B968CD3350EDA110E327EF065411CC9570E7C3501725AA12E17E64206BEEB73B8E8A82E43088E8D7AFD35DD5C8F7C4EA4724FE79032A2B4E1FE1BA6CF7A29AC86CEDC44849BBD39046E6FF90AE78F3A146F346AC1FB1233A983CAAC80F218A0140FD8AB476654DF560B95C967D43AB4AFE8039AA7188966F04C71CF548E4041E5BCDFBD86AF1347EE082AA7446C83125DBEFA44F5B9D73891AC89F4EBBEA04F9E8063830B7FE454EA2D7645D50FFD8A3AA418E354D8CA70282314ACC2FD020ED1432CCBF4AE04657E3C3DE2AEDF79C388310C7E3E5D27D2D2EC286086A8F7365C20AA8309B5B7BDA43FA459674C39C3C0B6B5F0EED83B54F21C7F21EFE1038142841F36656C9BA9AFB41D4B61B1BCE0F3385B8992979CB70F386093CCFC1C2E365A6BC31925434E5A646C79B3FB15577F81AED0E6E8065C66718E9DD4D8E40000000000000000000000000000080F161C222C343D00";
    verif_kats[0].PK = "3406C20EA187919F41CDDBF27F9C50A52B7EEED2870011EFF9EE10E8F69E0A39C794F3F7066E3CD63130D93950D0161F14CBA67DAE6D13A7DC8D9F439A6C626AD4005F3A48BA2E531C42E444E0C076496BC07DD0644D7096082258AA0D37F3D3D0D587E0064CDB9A505965691E27D295802D856B3295D4EA6562FB3247E343B1AE264E88A02B2777F92B64686F3F10C833A87FB693BA1F4DBE1812BEF2028BD37625D70CA9667320B8FBFB8C390BDD887A318E7AE9326BE4B457A612932C934E118ABC31A9C79D585AA4128E3559FF8790B96952C372697E96FAFF01E55168EC199E92A1360C3AC2196236561DC697A0599C072AEFD6A2683ABDC3C11557EB44B936465E15994D14C9B3F0E84EE72949CCFB9531F8CB75D79C9C2E68A1ACDB92C58A9C19241388C054345CE46CFC8AC2F1FF328639D09C071EB9E920F697943145B8FF45EDFBD8F5135929ED18091055CEE48E4776E87BBD62595E21990E72E5C09F48EB6F311773E523D395374AB1E0CC3D5B55F7EE22D2B189A882939CFE85694682685368E272DA8EAD2CFB972E4616FCD8143782C5C3A97F51CEFAC81387700C74D5D2E5B92CF762A1F327841AA117694ABA918FA29300C27DF3029EECC775EB2EA2E9EFA882A0EBA9E82C588DDF09FD4620E084756F5069BE893CFA1D8E0EC69962774E70D41F46F25F291C091BBAA447ACD24BDF5E7F0D6C50BCE69B79F51A4CA8FDD8343C49DE55EB3441E042404CB992803C2494D5512AA67A4BBBBBE765AD543C709A07EA71083EC4007E4828C58187C5FDCE680B34C902BD902A85E38C674B07D13E5BFC15CBD547867A3CC9A00D0DFC5219CBF4E82E7010B009493EE5672BE249DEBF2F4E91B5469F7CAAA5D5C69A080C8EF8394F06B8AC95FC8489A0A7BB21CAD3548BA524B609EEF7CE7C20DAB6C5B54B58307B416C3DB4D653A1446F25A8874A7B8B0AC6C2DBD175726849265103D455B1895213BA6C3D177CCD788145EAC23A65AFEF9CD75B0C2F0297420CDA46AAFCAAB92EE9955948A741BC3F60AD609A53BE44624520252957B2BA03113F6FEEFB690D0A7F5952FBB470F3F9075CF9EF0541A9B6BAA9DA6795BEDD8F41A27DF7F6C5855030354138E2077B4B2DDC570FDF0186DF23F077E1CF6EEF833D0E4CDA82709B69F9AC52E4D9254A7D0DDED46D64EF083C3585FA3A5B25D0323FDF17EABCBEEB64BA8513010494DF411045DCD48B1565697B0DD507450866E582BAE23C15010B6088806C254E6D81DFA7922F189F3A7559792F198A96916F96F78DB378541D02621D0EBB78C72D2A360E47EF09DDFBE1B2EC24C99C692E087D84C0BBBD8FF02275B51813624E97448C5FD294A2740D0775060A8F785630402DE3CE4357A655CB6DF2C534FEB3DAED1E1FF7C6161A0B0718DF0C2B3C228BB69D0D8828B876114B95621EDA905766E877DCE20756525A4C31FD84963974D984043B5A4CABFAF21297390A09FB6EC15867734065C7EF6B18AF9FB3596919820D21B766F5F2154E8BD3C74FD711C2F80F90431A44AE34997A9085765636D27CA3C3A7CABA01902D7554B0FC97180BF6547E97CBDD5E094CFF25206BAB14BF30C41EA76268996D4F011946387657B61E8715DC097DCDADE05A72712179F0A110E4203086C409090371BD175CCEC01DC33A7F4F20EF3448A1757E0C560BCD7747E6177346A8B8BB8F9FA7D04BE2D897BD3D5B5FE1231059BA5BFE40180A7F3ECECE7885B09970B692548C3D065BA17522151E0EEB32F3664C67D5164F92B48F3E167D71E11F3A822A2585BBE6395A9DD827933C31B7E43188830E5CF60381D6CC58DAB278AA0A5192F7CA4497704BF951000E3E786AD4AA651CD9E1650D0BBEE5B163287B44C1A918F6AE43C14E97A10E92F3F5F8596A97CC54094BFD618D72C433E4A7BC1ABBEA4406E5C5C8EF3FEC6F750CAF9654295FD26AFD89BE26B000B33C1F70DB955628AC16C0A25216942460A61A6807131EA5396ADE6716993F6D4D178B1E604DD078F2B488F784921467C3F93A4FFD2B9936F1C913F48B51EA64B64371EBC7B0F8A0ECA57FD0CCD614A130CBE5B9B2736CE5EA9652523AA2033DFF532F9FB94685456DB9C044C9DBFAED8B74CC7DED328737ED6D7CA13E55397699C8E0DE5DD7CA508EA4659C21A07968697BA3CCC7C9330CB7F8B95E7353D2B3374771709F364D82F3190134A27CD2A34D61869962F2403CE1F3218D9DA220B540F907E3AA578DFB60777A3109339CDB7304360E2754B3D07E132946C9DD795688A0704C75B10BFA36BC1306706353A1FD0BE5AE1560B7903FD411E49620D54DCC194D6E240FC87712C005D928B7A07C4F3337050D6060BA51EEC1D6FE0D7D73B39547E5F9331A6ADB3202EB2EF327F69C4A4AF35ABDE056475F4A4DF8728999D4D4BAA1650967269063285456D4CC8CE8C1F5B9E29E5305E387D34FB7259521E620D68DAB8532CFBF1021BBC8179F9225F38A0F04F19316F388DA2C4F6BF1C8F9A6343D890E4E4C71BA1EDB0B6D0B2FCCC559CC20AE06352C75E09A19A109BA1F1DC8D5CECA5D46EADA1AD47BD4F67FFCC40AC66DAF5B4DD15658B618631861EB6564BF13E9CEEB38225715E484983A706020875295D9BB289024EF61D116BFB84D72DD2D0F3C0373CF0605FE838B18E4A5D8DA5BD23D9E6E2B06E7044DB3D0774975FAFA8BFB6DCFDBE95EB5262FF93663A0A6F8A7B53BA1057E611FA1B3A3AF42741F291189CE1E2F628EDC1738767B0FEE93E66BD29FEB1C7CD9CE2D516CD9488FF33E9CE52198B05E2CD25020B37BA092F962B911864AEB5EE5E0037D9A5FB521EF99A1120B9A9F68A513C02E72794250333B68CC3A0AB9E473653D015CCAEA2B102B332B3B4BB95898440D6D290E73FF8F80EB40C2DCFCE9EBF64C574EFB9A1C3BBBC5AFA4D9F05F36BA6B44E66AF4959B79D706612CA98E689C56DB11AF684A004034FCFBD106BA1CA09D97D51BF20E2058FEE0E1A69B4A60B9834539AA94BA63EE1402CCF0D19B280109DC296CC2C40CF8441BE76C7DD2D17F3DE72B11C4AB7883FF352AC5EE4630D37BCD8D92291913F4B81021A094FE3DEF52824068C5FDCDE8EF26976B29DFAF51612837768A69CB3D06ACB1FFAA0B6F5FA0C5AE618D2156AB91F72697323A9D8BD3FE24A2B884B635CF933D2F80EB0DD48580ED87A30934AB5E7A5899299D366C09E7E3215935492E9356E3673E4DE1B29625FAD193BB53C0BC88BA55788A9970CC007288852661DCC161580FFFE307BF549F2721090C5B6424E9FE7852B8A76C6B06E9319B41720979D685669E95479467336CD68C06B48A6CB6916BE4D882D0C6371380F97F9AAE546AE520D843514E315146C7599DB5DF4D4BAA79EEF3EAF8C38EEA0DA201DDC5A954387C372FA1686F52C8F5CEBB9D54FF879D7339B5DE8BED40889DB44FBD9302BE8F0C20CB945389FE9B56770EE176D2999A9035DB69D9D13EA4E6F9CDCDFF55A5B6945604562915EC7C81D5D2B49E5B1750B01051E7532B8D644CADD714512948AA7F2D88CC5F154989A7D4221C67DB0852C02F6EC9A1EFC7CEAD302D871600C57CDD3EF134DF2EC0070EC7F8D1A80919045D1E630B426A941E15A0E1D6E258F47E2ABDCB9CA791F99885867CE36B6A49DA864A85A0C82B97959B";
    verif_kats[0].expected_RES = "277F05029232D41F8597688093A174585192D0CFBF99ADC0B2F2B2EFC34E61114B7C427A0E05C24FD7143FE66213225CD2F0D707B3D40F17BDBE0CA72D1EA0AA";

    verif_kats[1].MSG = "ca393154ce0e065793750cbb96156c74eb704ed0f2ac97c1131f250f550e1efab980c2cb146960dd7c0b562a1f412c6b2cbd203e1f048c73376590bd39d7a969";
    verif_kats[1].SIG = "8F5AD0CBB2C9E3165AFA169E719308B1474D6232C34BCAC63188945383B0422861F1B6A9F4B6F85AF18940C312D2D9C50C451D8A001F111D86A9C337F3A17AE062A46E6F23C28063A6B345CDCEDBA377821337E4E257037C3D4989C52E707DB4537B86A126AFB8022F3DF4C7CCDCED4D0CEF85FC7CFC7B0C8CF0CA48CEA1D7E9D14E2DE502AB67E3B36DD51AAC81DB8F8C4CEA10FC6ADADE94CBFA05CD962D701D80CD86D5F809BB3F5BC89D0982DAEE84743AC72A1B815C3007FD528BD5707A73F155ED1252A679390F02F0A88F4B6F9872544D381BE3D8B73D439D2E81179845F6BE1C5C688A87B27F88B680799E0F758EBBE360B90A0F4805019967FDF40D0F95F59CD2F5D4E471D2ED00718EFDE61F937E8537B6B25F8530C2635C1D11875D2C7800BA160473FD019CE8B20BD0CC842DD099FD5C7A815EF3DC8D0C89C1EC6BF5754CE3198141FF6F6A1CA29F8276A44339CDD4A0B61F16B31EA66E24D4AF47EE22AEBD4F97C53D2818D841C9A0638B03B016A0188BE513D7BE856FA563B8DC673EC7F3E711F7FE2C2B9F55D9BD372285633FB3013D709E0698637709F2233C0634D25B76654F6E17A2082F743B768B5E1540B0383831DB1811A8CA0F2991CC0112DEAA056D34949D0A503E0D69958EE9E921C7E47CD020F30ECA45CDAB485865DF4C20CEA5C671E0994BC2ECB740F86C9CF2443134F0E3570ACC318B217FC47D7F268D5F5BC8FEC5DE2726EA1563BE1963ACC7E9D702F2BF042C3F5919FAA19F1299F7E4C26E417DD7DF9AF86BB2FA82B125DCD3B35EBC3BE84D60D9E4472BC09B410A41DDE7B0950E0DDBE35F13A6ECCA3C1259785FF25A1B7199DFA371C57C46BA5C71D48CD3077318D65B07E9241077CC9BE7719A0574EC3758CD4DC38EA15322EFA6A96B022D14AC205222DF9C2FCF034AA66C390EEF568DCE0C8D93944EA4D27C725E475F63860AC4E56CC2D9F89B4F9242C90C74A93B16CAC076CC41B5952D367EE0D5205AB5C87FB74BA456B99A4A6DA5A733C2448E57B955464F4CFBE09CAEAC1B8CF7FD6F035B45809E1C24F5F1CE4A10EE493AFCB4FD8E7F2D32D50B400872C04643C2719EFB50CD184A91465F571D7FE770CA2CB21C4D2986EE5344944254F69A57B2BAC6B95475BD618CFFE7AD3B223E4BB1D9F70ABD7DFFC73F9E0A124FA16AD20A68A022C79A8164D74B68532A6986E9A97D09B4E03B50F170804666501AC6813420BFC352F839D49215C8CD9DA7BD7F7190FB12A4D117DE2AE664BDEE8B22F33EB1AA21826A754031593CE99E1A73498824E8167481AFA5660B3272354C69427C6F36FD0C0BF216F943C8FFFA8A132BDF7261676F69F07A3FC228C514FAA88BE3258C0DD0537190AD4DDC73B52BE3E1EBCFA3EFEABAB749FEC751C1DF235C6283FBEA4EAB9AC67FF9B3BA8BEF11D781B311B04DD7D41C44E2CBBF03F5BB6D983381E54EA52A986D8D535F3FD7D2FE063F097A7780BEACA3E2C65A02CBA89AFB09CFC6B8457F76864E6217FE49BE93F6C08EBAFD156BCEC061DEA3021C3E62B918A87A0C7EBC86FC3AF83E751892636AAF52C3C03A90CB944A36E976D1BD447AC88DCAFA847B7905B774856EF322BF1D7788962F21BD7BE047BDC7C5D78907483465FD80B081C14088C356C644299F732EC7D3182A66D32D53E2D8CE68BB8A355FE7B224EA3E12FA587E4B714F67B671A0B9E953779A1569FDCBCE8A638A0AB844A3E0AED8A664A784CE6D1B2CBE990035AA3AD943F0E90C6B580657C4FACEDC8998617075C81D506F24F342CDFE0E8390BF9F25F0E6DB9B4F5020317F534B5C7FD177E2ACD4DC8BFF8F785D596D4024EFAE44132EAF42A41BDC13FB648BC77EE98DD4F5B9432EA109027BFB7F8EBA68EF05D636EAD0999D8377E953F177CA98E2573FD7598D942F9620C17470F13C38BDF4B9CEE12DAA617ED4A0F38167C9F4663F5EB2A816B3DCE83C13E8D27939D2A5D75DF6484420DAC4D23059F21B89CC8960B798183F32C065DD3DFCDB187CEB90F6DD5671E8B5FA7BD9FB92E1854B309D1D2FE0F81203C868C10E57CE30E27A4B4E585911C85A95E5860F3DA3A7013B8BAC0E7C26FC7414F6F127F36B9F17329658D455DA9FF8D3E0716250E8E1CCFC495269A23A7E190F7364812AB076A56370EA32EDE67276EC3B6F245310FFE841721A1D7AD3FDA46B5D1B3869F58BF4EDC86EB182566EC063752AA1448AE664E5CF66B8EF172CEC6DF6F09B355A59DED9577AB2AB380B6C7A13B042E37515FF4728FEE4E3AC72535DE20183960F799BC7E9650C453DE6FDCD62CAC856CDC9EEFCED501FDCD23B81AF7122B096BD97678AA599C3C36347D07AFB76D15CC3F88FE1AD1919EF8C5AD329622730AF8C09D2864219BE7C4350A8170571EA365A7426D3AECAAE0498DEFF964A63D06C1C99BDD8650EFD758D30C541F4288576AFD7CE99D964C0117FCB2F444E7B6E9029FAA65DA3752B8EF6092BD3816DCFE3CD2B133EDF195C98883DC52B4F1387FAF505CCE8CEA2EFF17BC841179389F2F09B87849D55D516FF3DCDBA9575C3ABA2BD508ABC2772F7383A99FA57FA01416BF64A43A98D9BAAFCD2C488D2689F1C01E2CCEE0E4A5961D7FF0EE92D0CA4061BA021D9968FE0366743E90123F04521720725ADD43C46961DA9F571276711349A7B10D1DC3B2E0357EDB7B8C3D49DC35080EFD7A78915B8C0FEB0EA19D56E04DB89C55EDB1DF5B364566A5365A1078673E72957488ADB8FB37F508BD92BB3EE008FDAA9ABC4C55D73E8BBD8C26DC91606540FC69101F342196F395E45D423A84C29918D86D0F15B52E921C2BA97FE7E25D78CC05D6DF71DECD6D276D82C90595D75912E94148376DCFB80FBA067D30EB67FAD72AADEE53851272984D34F04AA944531E0F63DCFFC34158BDAFCB304C527EDE225C8EF9916744D7404F50416B28D4FBEE45C075965898720D766BDCA0C8ADDBCD10638B41E8063F94A061B946AD9F1DEFDCB1614774A086FCDD84FAFDE6D43D1BD291B174B78C80DFED56A4B0A4BD05F5DDFA5087E392C7FDF65EDCB3991AD4C6E93D424ABF21739868CC3783E3172640D2D6129FED1D3064485339C84A783DC1E97E09F80DFB34BB8B70C318C29189B9E32B614EFE0207FDD412416C8FE24D8558B4C85C3AE241E07FD54C02EA4EE6223375031FF300D73B75F729E42B17CCF8CAA1D9102DD32CDB57C0634E76083CD1C7D96F191242743652AFA9F45A84BD7DBD39B6A586A5C1958E802F1BC97E95CBDEE9E1CF5DB86DA648E462991DBAD2536177C8A5665A925036E604EDACD25F76829EE374AD21C2C03A0A6770774CBC43544FB38509A37F7985952206CC49EC25D7A45EF6F4094F098C96A11E9985C01F43DC19D159F5C86FFA78D19FC012CD800E305A4E940F142B1673C4FE692AA33A6491DD9FB8ACA7B46D15ADC1741584F1CEA86F465229C579E58A4515B02E51E2F8118A3D079892265B5042D438EE58D7223C23B5F52D27FEAF6BD7C05B55345092D104812628D49E9304151509729D38604A063B938CB3FEDC894D348024200320845F5156756463343B283BA40BE31F840FCA1BA1863F2E93CC00C1A83E666DD246503EA5D8152EE1CF6BE492559C360EC2743487FE739E570D8C53BABEC5EFD2ADFDE441980D82E6FABC3FFB29EC5DA8B36A459C7057DC031A556FBB746F6B5AC39857FE6E6D7EFB497BAB972D172E01404939A97048FA76084894EE22ED0491352141F7E98F19B00E92F88E332580DE46357A4FC45912EDAB48A9E4361AF83F4DE4122D6430F3D6DC5F219A657E7B566EBE52B1C68A7170C240AE806737BED4E0EC3D34A7B38445B8071E59766567592C7F9D4458E0924EBC96979595F15AEBB6A7BC1352C21872438D8AD2CC2DC476B196617924C97F85CD7C9561BEE75378DF9C697A935BD8EEDCF98CC5BDA7AFDD682500A84D5CB4758B48E3E3AAABA488798691A33E698C6A390306A9675B3E6440E9195968C29438B47E3182BE67E81409660F0B51F9A44D8730C070E4901D81907452F7C0B3D19B575727306857B933B736B69EAB2FA2F0403492CC08366F9DE393EBA62E48788CB3B5EF7BD04E4EFF91BE1DBA6E790A9073F9C4A80F336FB9B2A8E9FBE87533D4EE9BADE33B5357CA90D3258E87EB732F9D79D3C0728167F4E6E1858F42CCB7C52DE94DFEC8C277B0FC43EEB65DC7F01D074254C8F339F85265A578488A93DEF70735D0CC39D33794D3F60FD301FBEE3B2AB8E8182B36139DB3CCD3475D205FEE52E9E8C43BB845C1B213723CF2D53A96DB3BE71A65DC3B373126E16768FC9D5A575D1DDE62B79182AE2578AB0B56B042E27F23A574866BD52B08F0D6D836C57EF27D4EF3270DF82273B911A629C9F0FDB141D49F471D0B262D407912344309B1BEA660A6EDCE2A38C92245797DD99F64252348EE1ABD14A371695A9DCB3BE5854355AF8535948F87BB098AD116CDD982E492DAA5B07E8D9E51166CB9037FA00BEE764A92744B3659D3CDD3F69537ED7FEDC82440368A78F3C67700523BD17E55EF23AC5884AEC26D2879B6E79487B1CCC5AFB5A760B81C79988F62867BBBD5676F7581EB623996E0A06B8FD4F6BA6FC5ABCDB2D134F8C10EE7DB8EAEE278190B34D5CF3776D1E926AE206BF3C019CCE10F2ECFEF535EA4B0373BE58EFE1F7177EDE35195B6B43473F38D278F0147B008C4AE12F1E18D1B5E9307E390D0C549FFAD7237C98781093A9059436C5CE150EFA0DAB42FA0E16A4E1CDD82A6F06D97885D4B8C80508723D28AE9F222A195ACECE48375E62A4ABA428580006793A5DF6527F30D0F0377FEBE61577E272C26ABCEDAA40719862653960FDBCF2E9502B4213F41B41DB431E836BCC9DBABA679F2025584345B5192491BFEAA084AD7E4B2AF8B449EF59EC26C2A7C73317789F62E86C56F9FE775AD6C3E21EB6FC8F855872E0FCB71F6779F0EB35F56CA25A5A0DBD07B9656237220E940F0764DA242E27B59C8D7944F5DB71285885DB008962682D5EC3C0B01FB9BB016E1BA640E73E817DA3C76504AFFEF6EB9BF42E8B1DC14EEC14B151143438BCCD67556CF90329D59043CD68B6EEEA41A5231BF708DF78EF43D55E12EDEEA112008D72036B6AA95A94194EAA986F683A2957E48462A69A8D7B4040CBC84D3E06859ED205E910F5DAE8862E353816D3BB78D9933D731DAFBFF81541CF6089684979789642B449E456C7C3F31B0C9464A0CE3FB41EB809172CC00B37AB6EDE8BB0EB8B8B7BA62CB84C3ABF0A7EEE8CA0B92A4721D843D3F5E4F38CC8DA6F4B3299D08F98B07DE7F16F575B1A80EE019BC562E8962F94476E71C4BC10635BBB3FAC38F3419D7441B8546E08A588922304FB96DC14AEAE2BDBA660DCC0BF633DE7946755FCB437AAD79DE2A2164197A879DF640BFF025D0F6F39BDCB6C3C1E16618148B23DDB82AD0F1FCF2E1F122FC37DA0C280C31FDE267416BDD8976B847A1D336F424357C9FCE53AFAB9670BD2FB351615CECB6221D7EA2CDAB429CBEB3CC35FDFDE7E1A4946631AC85BFFE360BEE93CF35C81E3ACA768AD2248870DA2596D4144C593A2AB2764B4DD6E97ACFDF31693C26B07F8EC9AE2A58B6EA4AF4D0B3B9B5E8FA4DD62D9C826FBB7ACCB2BD2F1591525895EB1A2A02C822F528A0EA768924A80E4787E21EB763420A75A02CA2AFD6213C987473E7024DAED0B4CDC009C653643E6CDDEBE37CDEB525A1AFCD298884744BAD1C70D8CCA51D8B8D057EBB81D56CFAD43DC01F4706E72D62800AE43266D3DB9C8293EB8A17B4C969C4D6F8EEA47B9858DF55318DF4D7CE32990B5DB520CFDAF84A5DA0F0540F411954B74D8F9EFCF502219757D267FEC11F82B7092FDF6FE20123061F411FDC1DA2828D0CA0A26D7D5C63E28B9C81F9B10FF95E2B2EAF46F05B02F96B1A8D463908EAD0AE3035A102BAE93DD30E2B772A15482C13EF55F0A2F72724F392BB945DBCEE096121CD951627F8F801F9F23847FCFD6494B02C6488FCACC00B2C31A5CB8A26269C03635924DDF6B7C8A1DE3DF9B193546B9B8A88EFFA5427A10E4A8E4448AEBBFF4656F5C0F4E64177EF7A3CCE59B6073B5BF2A598A3617A66842BC86F298ACA86950A80908DF936761551BD13F405708F71B7370BE874D4C9ABE34D839387984D6606CFBB73206A98E997AFB220BE61EC0C18366508521B1EDA205CDB1F00CE26FF996F59864E29C6D999820D12BB03B3DF3DFA0EE1525E99C90DBEE55EC22F0042D0C15221CB5404993E29B54A3728383C7C89F49B106B22E9397E0CB55B903DFE90CA922C42EEAEBF0EA33633BDE99AA444E0CC75D57D4B12FFC8EB828DE807FE956E4EC7AF3383887398BB20FBEA3EF9A19B600A10F6758FFA22FD514D9BDBFC6B80A48F0E80110335CCFB78A14F5AB0C3520B9F7526E88732E22D300121B6568D5D9061F244059637C9FAFE0FE105F81BACEDAE9FB232A4A71D507273B3F8084AAEC01101C2C303783898DBBD20247A200000000000000000000000000000000000000000209141C2129343700";
    verif_kats[1].PK = "D7B1AE0B7AC9DEBF3236824CA48B49A5FF417C11FE65C667716FBAA44D3DD620F5EBDF9D49AF3B711F815E9BB80488C8F3106EC723E7CEE24F1408D73787A54AD9185B8A7E331F6085371C71C5A94A64B11AB9C2C05D1AB0AB8E2F6DE7A10E3562C28D10C563C57517688ECFCD7D2C5103511CEEB38C17DB88D256DFB1282A2A8D668543C2A5D44E01419F2FE79A9CF7708EEBADAE74956B0715E9FEC122CD98163DE1B961A79C343655957EB046E13CDF26C3E24D625F751D28E8B08BAAAAA2FD10D8071CFE63C875E129B290B2FD263D306D502AEDF01423A182DC1608B392283D0C5A11EA510048EC026E3D53A8F6124BA59929C7DB8AD898A6277218738C1FA2E51B338E7F2B7BBC45F5AB90A911C62608B663FD5DBD157BDF4C62CDDC3A82D8C07D70C896B37B56CC307905BE965B17EE996A1420044941F3FFBDCC6398E3AC716C78DC558DB07EC6AB6B2BAE75F2C8EE5A27BA0109E1993017D98B42933D19D9E0DE56D743E6CC681E2179A6972DB9EDC51902E6527A3A9D7C53B66AF3BA37D62684C0CE046798EC4CCE74224A1161E8F61AD01D44814E34ED69A77413414CCD597588964CD1D9824E50BB818928CDCE1FA35D470101EFD1664AB86A4C1FFCB2E51CDF2072BD8BDFBA7440BD9CB8643D5D8B1833B1771FF48DC532BE02D57181CBF38BCAAC0302E0B499DB4176B967973201E21B6E0E4D5ACCB65F1DF56E3D855F7AD2DB23CD0F838DAC241455A085BFE125FFB2526C3A71DB0EA64E756E0A5BCEB7992B10518AD366DBA6031AE43F4AC033129BA2A206ED17FECCA6747E5F350E0791DD0656125E682CFF2C0176F6A6BADFDAAEA474702BB1A60B4169F506977C693CB34DBA3010A0D26A5E6C287907E5CA1714A93890D9913D86EBC5900682CFAA0CF01573369AF40708F3CC83DF996CA12530B54958A288F58CF0D95C61D5E689ED2208E4A1AE20828D1098F894578E2C6FD1841A583954B037B7DB54DAFB11E6D8F38A7A091D777B36A29F90744C11D4DE7DFDD37E9E494E73C2920DCA5D8A377DA84148F0836C88D472FFD371402DE5A990D3E374F9478B834FCA975D261E79F9024DCD70DBDA745C776678C17B62353CD93A6380B849BE5680B679ACB0113C004A616D8E3208F89A52264319F973BA345E16AA40825D14D30FB179E8EDAF525AF8BAF56FBD44C97E0A3191C4D9A3DB9D4F9291BEC065988D82D39A5284F435CC2BBFE76367AC78E9768A12AC88F268157ACEFCC0FEA6BEF6E520A3603AFC090DC7D922D779B805AA38FB31FD95D656EF5DF3620122CA83DF5E83051CBCC2E6767A9005DF0D65DCD0863A3B6DDAA9357BF31D9E370A027458E687F6FB159935101ED576CC1A1965B51F1B46856C070F3EECA68D55DE610111BD831D34CAB4BBA7CBEA57065E27C2E2A075D2F301BF6B795CDD8C91A8610DC72E495A90419E58BACDAB419DE6CA5A06498E6EA382EC2CC284DEBF0AC7D52417CA1310484EE64C0C8385839D66A48821BC099BE9C267E0BDEBAAEDF2FED4C8D5C8FA38ADBD77B153991516C444B5D9F7FB01EA442B3F603F7285896C612B9332DDBA545B8342D9E553E7AB2C88A320F9206F9C72FE3CBFA15EC12541EED585484D9E7E0A97B44BFBFB66C48518BC31543C680A7D320424BB0A22697FE255E4787498F998812C712CF20DBE71750472C51D4AC501ABDDE8B90CA21476383E861721554A9E667360E030B02563E51973AE326BD3F8B9BED05272845B9CAED94188989624D70FFE5C6758A6BF6E225C641A3B71AED6F2844778C4BA844940544D8C8AB1D6556737E995EC517F66A60B616BA243E1739CB63443011A91E704210637807B72A993EECCB0C9719CD2FD3480FE45A4B329E7FDF51CC8FE9D136381A2DA3691AAABC604AF98465EF36FAB8C2C71CB9BD1C6D48BFFB072206903C6A41516212ABDD40206583ED0F66AED210023B19DAD522ADFE6E31586188566B7C64FDA5BC850691C75112FD5392CB18E5B1C2A0BC79A5FA757C5463F134980F2A203A93F759F3FD3AC4A17C71C5C6E428AB13DA82F3A52F45FEF60C7277EE256424542309C371B33CA9D1865E9F52D839FA9E578187B6D0C7390DB1715596ED24250AEB7968BBC9C5B77A73BC9B2C777E49B73F918D13BACF546942FF5070B760C1E624DB603DE558787F6BDB326B3C93165AEBE0B818A943FEB8B2DD72D8180917B739789B533FE057D3154159B0ABD67B60FF681E011E152BE6749F296E778461277F5AFE8BDF28AC56DAC78745545E3C20C8639BB76AAA76500E799078E59650FC82A0CB2B28A05DBF574CD9A50AB041D494A389D4DD779814A2B24ADF580880E95BC21DCCA392CA6CF7E9A50A3D80B5E6855A0426182489090BB82F1EA2150016B4B3EDD9FA3A2F8D85AD61AC2807BD814E5462545B82388A2CD33F310E316D4815F8812AC924FABDABE7E696E0FAFF17546F359430461053031D31BF20FBEF05A6EDFE9720E9BF2DCFE15D83A597B3BDC52714778176C3823364B383B61F5ADEEB770C3D1FE161407D697B6201D5F5B1121D034A6157E46F81342ABEE5D7BBB8977F6209219BA4B8DE936EC87054132CAC3FC65666199F48C20E2FD56B08D04CCD4CFECECE2BD1C65ADC9D0B8F26E5DD582845B761350A3A8E6179105B7906EA2DF4CC3C21402F0FD5ED1854A11CB59262819DF514CEC51C026A2AB9481AB229FE42B3A0494FCEC6C2F6AC160742254DAE4E4CEB4BCBD288108A71805EE27B994BC919BBCBFAE1E3436EBD6AAC2A56ACC37DA6D39B52266FD3A6B1331BFE9BDEDE19B6227575662CBD6DDC5049E205F30272C151BC0CC00E3A2EC4A0E012FCDDE6C51FC33A18C297F86AE61803B21346040099BE7B5F1527E9D648426F1A06D8F8F74DB968D439C04660B8B14EA5BFF205E273283FB1B40B47012E718C50C7E899533E591B54F8D0631181962EF810298B0C29414882E51B073B19BF1C49A893E6B541D61AA48E2EC909102C954FF63E81C40B61BEA01D642B869002D6D8BB1DD28090DB3CBCF1AF7FD0A17108C3842C12B4B55B741C28E303863F74B6A1998D18A7952CA6F1A6F83751A5550EB32A0F9218ACF9945CCB1181AEC15D750B74E6A6B170A6DFBFC7A09EA13089B6906CDDD285835D841C2F27F380FDA69A0679FF94715861146C9EA97A728E1FC7A7AC23FFCF8150F94DBD64F47BE44207903C64F2645DC7D4963CA94D0B97E395341C8EE2D52D015446F972415A5B651289274F57D55705B8152ED2948F8BFC84D7DBB127F30ACF4AE91C05C8D5C964992A4E6E8DE6B569F4E36C5B846A85544916DBBDFF6C9250C91B9523D5EDAC17505D6BEBBBC8111E89AB795298CBA5A0E25450EB73DCDEB643C051133408DA8F3D6B47C1AE23F1B010473AD0A2F62E63D05800BF9FB05DDB1040268A0D4F0EEA7AD172EF547A9685C4BA4AC0D719E607E96D4D20314153A366029A81AB826BD5235228AA2230C6C0DE15232F7DF8330536A5A156801ACC2F20BAD0DA972A9FB2B4566B48F648A9F870DE8181484DFE57530A8EB0E5C214C418224699824CAE98FBAFFADC7C9DDAF635ACB7C92B2113480FC110E1D43B6DDE1A755C4E11F197E7C8CFA38195774B65DB88FE7EFE0839C22617E0FE33139EFCE9342D2CE72616CDD58D0316C1694";
    verif_kats[1].expected_RES = "8F5AD0CBB2C9E3165AFA169E719308B1474D6232C34BCAC63188945383B0422861F1B6A9F4B6F85AF18940C312D2D9C50C451D8A001F111D86A9C337F3A17AE0";
    
    verif_kats[2].MSG = "9433ddf6e491cbf5cb03720b542e432f868bc7b5a0bbafd914f210c3a9d145953c6532b8212660ff219cb0bd283c6c25501aee58ef4201916e7671f92b759f21";
    verif_kats[2].SIG = "0BA12A7496E9F3553D01AF2901CF4C423AA6F539B0FBEC61D9FDBAB11EB977ABCD3A191BB7D8869848F0736B89CC1221575C114F0E51B4E636178271044092579D793D39EE62A3F6DA6BB7F406BEC5DBC83E6E825990DD833BD2C8B040D084B52D9576FC6D950E9AFE96E861BCF6307EBEB51B13A6B5C1F76F2197515C5A2018E6D7EB45D7900CFC3F70D29891DA1E121FD45077C3A2F87E90E9C98F7F4893C8DD423D54B91BB25C7EEFB29198B09A84003CB375C5B164C670B4331949111102A68075747BA6AFEA02760BAD029D2AD02230C83296F35B893E46F47AA8782421E98EC0A99B4683A356A5BFA780AA6A6F9446A0E185EC98AFE12D15D5C74FE8BAA653BB55CDC37565463BD672BE195B6BE6EBED1670B691854B539F5F1442BB24132558D01BDAC6830C7C7320B576DA796BC25D1A00A96834E3A8B014BFC14F30BBFD27F9EEAB2168EB4E692D03A189E3900C9EFA98ED66E4B9202535CD29EB84859AF15AD66D3CFCB7FB8D6AEA19D9BAD2D4C28ED33B868376DD0CDB9A5531F5AA556D691E5774536698670A1470960CD3A2AA0FFA7628C23EF96A6786EC91A050426F54B36FF846E1C811631861BB32F49147B07C78AEB18991A3E5FBF8C7F92F8530194CFE1B615FFFDE26F3F727E5B20199F8B577888AE112F84C9A0189DA0D6B89636DBF696BA1CF16FFBBE1580BC0952903EF69ED922640E6D0E7B3ECF816F39D06FE6FE8EC98D31D305B7CA362C011E3B6FA1599C83B36CB60F88C6EBF1FC3A34DF524DF3C7FC60AF3ABF4BBFED3DC35964C2280E2EB65689B4DEF57E913985499EDAD84A4C66FC4129ECD660D12270A8D00C04F57C4C786190B69A88260E5D2B5DE1E2F5A39F077F57D5ADC8AE7B7536F321B7A91971873EA53761C97E94CB0B43C12BBE7989A844469CC3BCA46869879FC577CA7A7981A18620AEBE29647EBB6015654DB05A678B9F58643CE0034052800F8B48D564DA7C3425E58F2A82612323BD31CA7286A6A0F9C80A2C3D593F95CF5E5A4F16241AD89E6A2ABBCB3DDD1DE59DD0024A827E66C2AFFBFF50CDA7D4B9E5921923892715115B6AD7741F3DFB87FC57DD17028270822EC9114938457737584F2D57FACE64E9D9F8575855F98C8D49A10D5772E696486B01B44CD6A383A255D94FD07ED2CEB7D933ED7ADD6BC274A477669179B9B188E828A9457E5A1B3E38CDB6719C34506C48DEF82D58873CB6E6A76AC5883A9EAAB520B6305642081677F3A1EC2AB5C35488739BE6541A226114C6BB4647A3ADD06DBD66B1ACD2D775ACC78F89B70110A0E06420E4C420971D2ADC5F5297A5318DAD009FE042674A186DE1B4CE0B1C1527118BEEFE987195954EBD57B93A27A281B3FB2B800295A2185636D99DD6260290863514346A41125DCCCE0511778A6AD6EF93987A32F6010A114C8AF50E56D9B1F223FAA45886A3F4B1D06BFE96CC3B728CB8A781D465B9957F19B075E3B68E83F6909EC2DFED2728ACE7495BCA341B930208448CEB4CA921BCECF94FDC84E1BBF56AB528D8696A05CFFDC3B716E8C36E244F69FFC757FE25C2AFACA223AA20DA115BAC88BE9204F53E2968D3807935039D36EBD6391ABD82FE364AD41CDB4927E18128BBBE2C014166830CD476DDCAD141E41AD5CFF8D88939A157C65983EB76BFBA253CB94A17B8C07BB2388DD3C0F9FB2DF3BCF25B60A97AD2A5DF7D4CAE26C91652DD6A52A3C2656C6B5FF19271B93DFF1026E8069DFD626A97C7FC0C5DF4CD3EA029E1CE510EAB1980DCA4957936FD6D9FAD099FA6A898E270ECB5FD1D5C1BBC5A4803BF18B23532793CA25850660965386EB3C281CDF512DD64994930CE2C81731B09710935379D210A8E6BDF921CF56BC6C90A32E1E788723C1CF9D9416A478814CDA035CFB5A11EAEE261B8CC5131F818D39AD7C0BB0A9571BF5DF089F1D4ADAE989E71F75610E9B5EDF067744E6632A306AF0AF5B3FEFDD02E170619A7EF50585C44697FC7443A3E8832A2307CC8897A114D6C2E8E51350785993695952F8DFA78F2E8425E3751858C4FB763F87C032A35B459321325E6AEABCCFE96B4766B361E7C853C75931DB88887CDA86D7DBFE512637F7B0623B5F83DCB970D16E549D1DDFDB8D013272AFC331169DF5EF0F8861434828213F26429D47B448BA3AEF1B484165367B7C0AF999825D56FFCA6E6311787D1B416839EA96CF7A601D829476E50A2419B89157E1FEA7708CEDFBEE5997DD61702CD05AC3A9F91BABAFEEB17FCD5FF58D2665D99E735F8AB4DCF5F4C3347AEDE1601FA24A60CE8A90C5E371E1D118E1FDF68B5B57CF141C339C1F63DF5D6EF0789029052308243737C395FCBC1E91CD092B40B28AEEFD915294CBBE8855BE49182B723BDFCA0C824C1F7F80FFA1CC7725B4595A63BA93198B07257FD95FA173FDA8588E30B30A06447669D480F8BFBADD6945470513DEC3DAAC839BF674802B3CD467C6B33F916B708E9D200FF87C5A887E94031EBBC19E0E98495C5302C181A165B0959A20D4138101F0B420BDD1F54B867BA2618A341CB3E473EAEB23FDDBD2253A507C9DF628D91E70531193903C162504BB66A6CB291D29C6EEB478211C77B88696995B3095C090E6F690CF9277909488A39CF0BD72FBF44E1DC38E7BB333367494FD2C0ECAEC91B0355FE98D940C1F00DDC96E6E9AF830E4528E637A058FBE9244CFEB52C23598383FB9BC53BA252E656B9DA1B62C730257A4C737C7690C97EF7A3419F80EC7E794086BC4942096737CFB5E350972181CCA3052605FDC5CCC3F4405244CC299D88BAD0B559B5E5898F1650F51747D178F96A467908FD431BE4C07C920A0EC3480035D7417272FC8D83A60BEC31735805C565C306E5C706428DFA3E3A34A04608738B63796FA74CBCBCE7D472B1CEC8B9A19793F0E29BC226624EC93D9C6A83173DA50297398312B244E2C84387E3BFFD68801954D839D7E6598B28661DF19CAAA0E447059EB15F65E36A3BA4F8BCCD923A5FBECB0524FB2507A469D33AD51A7362F48F6A38056CE75A8E6B946D30620EFEDF3BD83E0CAC8B45C162369C4C9300BA4CCE9965BE940D1386C9913E981F6FF06F2DF3BF2867AA24A008EAD24479DC324E591772D6B72DBAC90BCAB11D9E16001E565A09D36F12FA81A7DB79CED92668D3248EB391FF123FC5C7EE1C7FD5BF7266D225DCF676B1F3B2DA7B4848DB50B2ABC75676551D0236614A3DA5F731A4F8693351716EB5CF95ADB76A5AFF6B7134ED9A569A3D575B0C6589BB22E48075F6297B39C683D50288F53F5B461FBA9A9802CAFAEBDD84359E599B3F54C71B631445CED6AA90AF3F61C35991E54F96411B66892FC609A9E8D58218D4DBFDED5B91E8EE5D92CB1C22E363FEFCC1E4922C2E094597E2AF3C4D771E562C7CE221A8708F39AFD608695E443AA8404E3363C429D4616D7634BEDE5EEE106B6A3E6928AADF44997ADE04FDA077353A6C057FE8E9BEF3BD4688A798B5A2DF7C491BF0C665D630751219C0762EE102D70C5451FD3AD50A820BD9326CC4D046A80A1CD3BCAD8AD6A246110CCAA71B581EB140A60853A796252EF29B19913D8A8E78FE66616FEBC72CB0967376A4553EEB9085FA12890EAABB251B7B8CB65C859602E4E19FF42AFD64141CE9092E4DDD937DA5D6C0C3301DEAD1E560E6154527819D59C915571999363BBE9F209D2217E17379F03114236159D2B1B7165B5503A93FEF37F3193080306B401B6D0D2084794FF19FF08D181CF8535D6545B5E30AF2D6E5356FA158EC19061719D313A8971EB85205C7923F79FA1B31B095EDEC9C8DA853FB3D84AE288762F20DD923B8C1783C567ED82E9B016048026D86C80DFD50FD3A2938CFF6DC8F6DF69DA25A4676C40596871831C59672F84F255B6A78EEBC67629418D883A88828DC9397CEC0A6201E6F574A57826634DAF722D2C76AB546565922041226CBFCCAA8128766F2AEE002A52BBEC2452B8143EBAFBE9F04B72BA1B085449C742FC42413C83952BB51A6749462D55719000B88BD9E2502D5B5EC77D2A6B11051B4F1A89C68E2D8DEA4D82CB23A29158DCFDE17CC42CAB7666A19378085EB619417BBFAB148F3A4144D9C7A7727388952B9B74472EEDF9555C88981653DC91FCB1D9AADDD626CCAF63D3B63C6F95600B7FD7AB16C95BDF5459436A643118497002DA57BAFDE6C7A074729E444B42A53F68E9C81895B9F0750AD499F73E47C519AE70F7F01759F423BCBEEEAB932FF4E4A17C140F3A81390EF4FBC3DCDAC05690DE3F219B7FECC900EB8EB7F268B3CF18E2981D07F7CCA4BEAECE2CFAC998435223608F06B3A1CD8474975BE376C99D122A51AC62F20D16F177BDA0FC507C0FBADA3E303E6E2202573B22F621F020E34ED6F48D1089FE65C60480108FA426D1DA85B9DE006B40773D5B043FDCC10F9A1F60CF6D501D69A3D1AE3250E1782A8A05E4B3A73D901EB8FBA9151631756B3F4622C04F77111A294B2372F921B28B22CEC8F31C95B5C09C0FC37300E012142264EFAA7BE248887678D4854626C6BAEAFA76FDEE65DCE6FC429B35EEB79FA26C71EA8E83A7732A65C854CD2B6FF50150323A507934F5D18604D73B5CF329C21E53764E5A7D6F47998831497F4217FF9EDF66BBF182EE607BE0CF6DC6981A2E151F460C2A43655CBB5C74A0C5175CB9C2491277A483915F9DB5FC435B88B436E195FD9B4D8C9F1998246F463431079F4A377666472209F6AD8EA2C69571528C3045FF0A49AC9797C7B5E7EAA7151C117333B335793E7696079A4E9BA2AF66FD1AABFA7DA1DDCA5B3CB010F8DF7A6EC1EE1CEE52BBB6D4E607D8161316353B71C0E280B9E055026CE0F70BBA372F2459360CCC767156BEFD99C3B2C5CDDD1E1347F839FF2F8AFAE7AA54A1438DED82E001D61D0B267303E2BA4C6CB6F2B449762D46710A56B1E22F3127F860E578494C48469245F2FCBB0E43AECF8318571253E2BDFDC9DEE1F35B2393F5AD2CA338806A0DF2B735F9349D7A9856C944C6D1ECE3795A26B3605693C69EDD58C9EFE6258A7402A94DF44B13329A419B0341FA1D5266B21FF9FDAAF8B6A5C933DECF3D9D84121C4978A2C02E249C97F45770D2F04BE37B0F8632F841AD0811CD276703AF765F4DEE1E5E89E0EF598760BC70AD3BFF43A216EE748885733F446BAA3E8A966DBE3DC58E318FEB2B0FF79C6533C8467CA0F2B42E7462C70E335C0BEEC5839D5CE84AF91417E88518A2D76C3E3DAFCDFCDC07FDBC5E9CF5CB11B4B22DE91D55CF576728B6DDE42039B8DE95B4FEB4372C423967FC77349F7F686C1EDD8FD8BB6ADE0DB5440D20B2133E1D5176F0E4B9117C44442DF6724E80DFF1D697C4ADA4B0A119695AF69AB9DC4EDDCF34D7210C3DA05D36941260B7136C67BF937FB01A0550C23B9DFA1A9E49785D994F22C3EE2BAE42749F2A2BFC7BC5A7674908B142CFF56F8335DA4958CA2CB61C7A14A64E90EB9B162E4E51B8976B237A5A1E077192B8078893BAAD319143D9E696C8763EB5A1BB3D32B547131138D3E6867A98DE044E374E9F299D1737E0366BC2F81FE33E0B1D3E3C1EFDF48F160738C20E6E9937BA1D39146B1B151FD668D3298CD88C0F9E480ED322936B1A84EF2C5C13F2682AF21F8896B897A66B4F2D045BB5C8CE2C1BC5DA9172FCE33346184B4BA27DAA96AD79823BE76EE26735A30E73EAFE17B5708C4AD770D3CE0014BBC7A00D58328431EAC8899A1A36B9DFD11656BD06E97529838CF2697B897D2AECB1C704CF55CA8EF0F38941278F2AE6DD88651D9BEBD81763023A88FF17C8C67407BC3A07E1CCB8DB1CAC81F8743A8D5CD787AFACD998DC43B39E11734A36BE855BBC48E1CDF7D8CB93D1646795E4E433A1CE44CB52439EA62FD0C80D5EA9072F51F454A1C1E252EEECD9B3E081FBEDADB6E9EEB0F110DDDFEDFCC0AD5E9D57889C24E574AD3C5A7BE19182454C0A1199F0C8D3ADB92A86F109B069A9BA74B8060A887E34AC58E0419108A945BD93DE9CCCFE84C0E8661BD75B4D3C059B7B5B6A63F6AF5E2AD6B4C7711FF6F57C582A871025B1592E32010D2E2B99FFA7C6BB0635D158914C792BA71E2C23ABAA62C1937A33C9B1741C3EF222D719689BE9AFB2D378F1DF29D97087DDCBAFA9B5107CD7B816FBDB9284905226B9F1F0F3F18BF4A93A2B826980CFBDD97C1CC758B1DA0964E51F899FDF99541D8F75DD5942A2672E5C1503CA3114F0E7F5823DBA847829A04DF923F16A5408961FA60AF2E84749E05D7F8567104F2EB3447736118D67C64B92DDE6DE87AD6DA0506ECECB5E0DC885664046B86A5D1320B82CE91D788C099316634F8FCAA94E8EE340EC13AABF189DAC6F2C7D4DC66C44DBD0897B19ED072B009DF3C388878A492E956BBE31D85CB2F7EA7F4E7E39838391DE84AEF020C60D04753E8724EF2B695ECFDF0B3D48909BD9EF23376B6D7AAAAC042B2F4D5464797E98FD0D3C3F5AC01A4A5766718F020B15216B7275A3C3DE35546B829697B30000000000000000000000000000000000000000030A111B2026303700";
    verif_kats[2].PK = "58E3563D36F5D0492030B6E5AA317FD727165ED2F494FF5EE45F7E395045C87E4B5709DFA6E7688B11B81F70BA940DFE52729C62AC9C8D56B0A93D2D2EBF4347144EFBFCAE4BF801CFB1BB6570A8A58C27602F44DE8399E1EF6281B84DB2614F4DE383BCF4573F411FF97CA729BD3503FB2F91F5F778581E89A8A44E3C3C3A86893E78F991B7A7FDADBA06C938A8FFB66F58CE9B584FC5DA89190BA94E896784834914A4240BD8143E1A12BB78036168B09D1E4BD274FEB8084EAF2913617D2A1C6BE16B54224C552B7D410A831941EB25AB9ADEF774A1F73FCF1436D428E051C23B2C7B08CA788B5A70768FE2B6B202139177A153867A236A9FC9CEA37F47FB7E2FF30972DE89C0850DD7B38AC0F855BBE607FDCEC0E4A32E7928450EB1A571357AB0E137830379F9BC7AB2D8D25C3C59E56229A4DFB1B28BD9B7D8A0B5FFECFBADF3D24EE4E15CBF34D6E771AEE04CB3EF866083FAE94A7BA0853AF896B1438FFA79079DBA05ED1326479B79EF1B770057907CE068B3A62170936F42DEA21E596710A0975BEBB86D605A8A1A4612E47F9E60678602080C57D07451D6F207DAC1D55444892DFC4783FD0ED05DC61054D1E5E234D11AE559C35EAA3A5F6F2EAC9F908600FF2229F188B3C7C3488C88C891A0016198F6DDC951DEC5BA79D217A7779D18938536B8A049A8E418E1A73B77490A8A11A7FC28F100D3F706EB490AC59E38D39F30BF632B458F4CEF494D5132D6C74864737D05AB0AC85C34C91A19E4BC065EFE5BB4F27718D9FFA0431E5619F447CB8C92111EA5AD8104C57C47E5BA02985D0DFDEB9BC9A6FACAAF57F4BE0BA680BF83308306BA43838F7EB9A8ED5F1384134902DE002705100E6785B2DA943ED591CAD0A085A850838E10AE9889FFC1CD2941E1899E1A26CA56CB7480D260B217798056D35EA62BD55F159CF0FC363A4F325235ACC231BCAE18E89EB70A6970B2EC08DB004961FE951F8ED294D7D68CA6DB402325D054A47D17FF5B38734298B99278273021F165817E7805D581A0B9E40D507CC89D543F7A1B718820B1F8414AD6946B1AF7BC3AC1A520312240C0B499CF6B2742508356F9C366980BB1894D343E1BB24F06EB81CCCF5CAD59158FFD2C0D5E0019A839EF8AAF32292C33E32F6454BC03F7CE05D157BD875210A4276EE7C828291BD5AD5D545AE4711FF0C1332AFC7D716D104344E88BE87124ABD94216405A370AD8097D80879DDE60CB1F70B8F2230CD81D719EBF1C5C1D6EE965A85CB8C9982CF1625BC69B0C89D5D4207AD037DB73A929F024DDCC2306CAFBA0FF819CA596EA988A366901172C153D7D2A467FA1AC7E738F3335C1A2008181A8EF3064227FE7E72DACF26BB28816BBECFB8224167224BD37C5B55BCBA256C9CBE8B18FF4C36EE6A1EF091A714416E91DB1D638592D0FAD1DA51085D36D12B1255884B849B2B6C661A9FACBBBD67EEE7BF27CEF998FEC1CBA2E5EBD5361B429D509EBFC6CB2DDEC67B6DC69884A342D4A6C6D8001E9652A1486B5360A17BBF3A47DE94D1A32A5E2602FAF1A41B5908F67E9832382E87C9D432A3B8B6E230A58EA733F980488491E7043F327160FCB6D34383FEE41FE7DB76D5BA72B3DF23034E648E8ADAF8D53E1F63403A62CAF6AB88CDBDDEC39E9AA4233E3D335DC890DB9454CDFDED997B292562B5B001451729C833627E9FAC08097FDBB64464CE6B4C0D33FE64987373951F2E3E19E7CE119A82C2529C244BA56C7BA3C703CD7C940759403829A505A635B4401AAC9A8A9C76EB375F6069D6C3FB6511E20F1E9F1B40EC3CD47CB90B638329F17E1A3D9CC45769AE2E6CFD9284C11F4B0892BEA676F9B09CAA8E83CE7B7648546FBA7E7A8B9580ECCEA43FE330A0F1520F5933164F524CA22EBA3889A51D184885E515CEF8B35E65DB4DFD90D8D4FA1FBD0F7F0936E55643905AC144175A27F189865C011D8570E2A57392A521C6C38DD7CE0D3FB5FB4C34FDA41645E5BB32DF8100507B8C0B33846D12C5878D5AA05B86E4D83718B5158E67B4D8CEAFEAAD3760599C63A0594B64E21DE4C1734AFC875005B798550F02D1203D94202AF189F140D3729733C276DBD47DBCC0B427CC113A38382E4044B74333D6EFE559FA327F9EB5DA8CFAA99B882EE97280E7A909E4B23A0D35CA8164440B71699D82623BD542ACF364C6D74E4D8D79A0C293629474B5D8A05D3408423A17B9045E9A3A6245D4F123DA541FB8FC8C5BFDC3E6BC508B823DB3EA81D1529558416E720346DEC470E5A7FDF7720893EC139DF5B8A7664ABA3FDE76AEEC0EED445850B5FE0F81FB3D0CB9BFC1432EF66FB8960E4601B50FCF176AAB7AE4C0E9328CBD5ADB4D8DD89DB72B0221382D96C04A8F511659D62FB268D781EB68962D2167806C73916CD66DF16E9CB7A1C25C794953FC3C87326AC3195E6285FE5076C35A56F24E7583E985D51F8EE8CF24AB0E78F2873E426C20B94D15A1E178F22D96C4EC22E90EB07EC066CE4A19BDCD66D03CAC9DD906D9D85C630A7E10F118D83DC7618AFECF90F3CD32D265253A05FEACD7DA610FC868BCF54F0053BB7625CE2E2C35C8A24BC8F3DC294F60DF8F345ACF03B2D8BE69B36E51B49492E8891FC09787527B3BEB02E6B2B69158448AE4507FBED5C3FEB923854656B642CBE0176DEE52B92EAF411B5E1480738476037D52D7AC9C04D909EB7AF11D98BFC66DFFE81F19CE1AAF2E3C646679B834CE0030A6E3AC7BE93027D2D7347B9165F9DEB26CD54F33A90A3AD5FFC88044202208C3D1C97B9668542D6F1DC4E1FD2DB6489392E9ED43FA989E5CCD6CC63E357D516167691AF5558541513B38D8DA32D19133EDF12E1D161C5873BB423B4E52D6B34E97875186D0DF7BB4EF4D05023B19274FB1DF47631F6282A45FDA95A07F8D5B0B0F814AE31CF30947FFA65D940C88CC191B3DD031897F8647D0F8D68C2FB79050F90EDA905673B206E6BDC844875101AED46513041695E9EF151B06AF764BBCCA82B0C93B9D26AB96877B49C9368C972E5D42E2CD41B3F7AB17F8F0B3EB1D0C284C699D9F5523D6C5E2F1E33747E49EB675CCF1B68D2CCDF4C7CAFBD6B1254C141001BDA1E8A9FF6F05C8B914182BC4348655D69D7DE203ABB70242AD8851369AF610CAC22E62A9B300F53ED948BF17D811B6C6B65F2E858E645F95A7F2DD7A9A6D6C2D627BDDA4C852C2AF523F9D03109335639009697FF25A1C67E3100083BD6A741A5B4C8D5567A85820E3D9CC6A7F03A1B7C902C75EF1DC49566A0E3A12671097F086CA024E61DE92F15303B0D6613EDF5FF80A5AF17FE2613437263899D8F66DD19B34A7887B72F416B8DFF7498EE37590DE4B1AA099E9AFE8B78D139238AB3473B60BCC70616F6ADEA0CE912C640D4672C4D68F2DB405ADB6643D7C82EF4F4C95DCE932DC8C96C870B1B7C0B91CF5150EEEBE6973068A3E60C5DE142C96A2DF5495E1CC3B3823608116D0838A5DA3A8AEB40887C08E58A62EA753FA3DDD0BB615646CC2A5B185C7B55A7DDFA9704C4FA0A74A2B1BD579C24AD9110B103A6042DC329CBFC728152533A41C3DD19C7F07F5DE5C863C97DA162E01FAB8E70DC91996897C68A173610B61558F298EF0A540BD762754DABD89B89334A2F95A9861879E0D23DFCA4DB8F04DB6A7E6A3D67";
    verif_kats[2].expected_RES = "0BA12A7496E9F3553D01AF2901CF4C423AA6F539B0FBEC61D9FDBAB11EB977ABCD3A191BB7D8869848F0736B89CC1221575C114F0E51B4E63617827104409257";

    // Iterate through KATs and validate
    foreach (verif_kats[i]) begin
      parse_hex_to_array(verif_kats[i].MSG, kat_MSG);
      parse_hex_to_array(verif_kats[i].SIG, kat_SIG);
      parse_hex_to_array(verif_kats[i].PK, kat_PK);
      parse_hex_to_array(verif_kats[i].expected_RES, VERIFY_RES);

      `uvm_info("KAT", $sformatf("Running verification KAT %0d", i), UVM_LOW);

      // Wait for ready flag in MLDSA_STATUS
      ready = 0;
      while (!ready) begin
        reg_model.MLDSA_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", "Failed to read MLDSA_STATUS");
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("MLDSA_STATUS: %h", data), UVM_HIGH);
        end
        ready = data[0];
      end

      // Writing the PK into the MLDSA_PUBKEY register array
      for (int j = 0; j < reg_model.MLDSA_PUBKEY.m_mem.get_size(); j++) begin
        reg_model.MLDSA_PUBKEY.m_mem.write(status, j, kat_PK[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
            `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_PUBKEY[%0d]", j));
        end else begin
            `uvm_info("REG_WRITE", $sformatf("MLDSA_PUBKEY[%0d] written with %0h", j, kat_PK[j]), UVM_LOW);
        end
      end

      // Write MSG to MLDSA_MSG registers
      foreach (reg_model.MLDSA_MSG[j]) begin
        reg_model.MLDSA_MSG[j].write(status, kat_MSG[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLDSA_MSG[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLDSA_MSG[%0d]: %h", j, kat_MSG[j]), UVM_LOW);
        end
      end

      // Writing the SIGNATURE into the MLDSA_SIGNATURE register array
      for (int j = 0; j < reg_model.MLDSA_SIGNATURE.m_mem.get_size(); j++) begin
        reg_model.MLDSA_SIGNATURE.m_mem.write(status, j, kat_SIG[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
            `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_SIGNATURE[%0d]", j));
        end else begin
            `uvm_info("REG_WRITE", $sformatf("MLDSA_SIGNATURE[%0d] written with %0h", j, kat_SIG[j]), UVM_LOW);
        end
      end
      
      data = 'h0000_0003; // Perform verification operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h", data), UVM_LOW);
      end

      valid = 0;
      while(!valid) begin
        reg_model.MLDSA_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLDSA_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLDSA_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end

      // Reading MLDSA_VERIFY_RES register
      foreach (reg_model.MLDSA_VERIFY_RES[j]) begin
        reg_model.MLDSA_VERIFY_RES[j].read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLDSA_VERIFY_RES[%0d]", j));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLDSA_VERIFY_RES[%0d]: %0h", j, data), UVM_LOW);
        end

        if (data !== VERIFY_RES[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("VERIFY_RES mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, VERIFY_RES[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("VERIFY_RES match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end

      
      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end


    `uvm_info("KAT", $sformatf("verif KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



