typedef uvm_sequencer#(ntt_txn) ntt_sequencer;