//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef struct {
  string MSG;         // Input MSG
  string SIG;         // Input SIG
  string PK;         // Input PK
  string expected_RES;  // Expected Signature
} verif_kat_t;

class ML_DSA_verif_KATs_sequence extends mldsa_bench_sequence_base;

  `uvm_object_utils(ML_DSA_verif_KATs_sequence);

    
    // KAT arrays
  verif_kat_t verif_kats[];
  bit [31:0] kat_MSG [];
  bit [31:0] kat_SIG [];
  bit [31:0] kat_PK [];
  bit [31:0] VERIFY_RES [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    verif_kats = new[3];
    kat_MSG = new[16];
    kat_SIG = new[1157];
    kat_PK = new[648];
    VERIFY_RES = new[16];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // signing KATs
    verif_kats[0].MSG = "afbdf91c942b5eb73b7cc474e53c05213fa41e7a2a826c58812f3065e7a289a6bee9169d145d9c81fbab6bbf7cb65e26d31d734e755d7abab5db81ed9290fb80";
    verif_kats[0].SIG = "89E8DA09EDD3600C15A06D5B5CBCA92CADF08F4313D0C0E2B23E24B329EEBD1D81DE6DEAE3F36797A494BA2121E0A274C3988770902E2CB325B79FD1C6ED2197A6386D50174548C5EAC449A1166F864DCC6A72C69CE883B783496A8FB7D7CAC3114996337082E3D45913F54151184FAF4CC4A45E71055E82E1F07279006278D00F427C1385800609418D46A6AC9EFC88E65C6532F2951B4C54A3EBAC4ABD047E9DBAD4ACBF9F1B67F53CDAE7C95D59CDE964C7F1644B2F2A2F2F3E1F8AEAEFE0FE7F6BF620E04ECFD0C6409FABFC71055B31BFC124441C388DF7B277DFF16EAAAD5985807DA361007E3163646F44541A623271B24ADB351CF68BAC7EBECF63B6C0ADDCF80EE0440BD7946E95F188C2DEC36D329524DC1B46738FB3FF0DA06FD3944248422394569D3CFA33E65CAB3E8C61DA6256DD396995BDEB151A5B7CDF429914F35FFA6B796807D70426715AF96B379DAE930D51A0717817CBDA0EF43F0EA2BEDE04D9FD2C72870F2B812818333C5EA491C344F4D359EFFC91984809A74E431DFEB05EFA1BA66924E4DEBA91E970A3ACBB2B34E272092E18C4FF4CCB7302C0067CE923C68C233AAE99B7090B7038CEFA82AB19A34B94D21FC70A8AEDBF26C8F2A4A4B74126E3A5E488579D639ED3881308E25143C2DA100395CC9F34CBFBE6770AE3D48C52AA2B9E1E1FAE2F6518E1BA8FEE95A029F72385FCBF1E1FE3E3AC96EDAF345104480F4CB407241B52AD07D896F73A12DD5123402E7F7D3E1B6363003B2388A351707836936A99FC26E5616583C101AB886C4A4B519145509DEDFD6C0BB3764B0BB3DF86DBF87437232C63881A74111058A5A415CB0708A20DC180391813D77D9F9F6E4ECB51771C101B2BE44701676D492E5318E995E6A8904657958A8AD1B11D6DEBA66DBD20D2884E23818609571EE5908698123B2043D813F1C61C6C758CBF58EEA1D3D3C7A01FEDE5E782BCF5DDB9A1CDA755EC0606D4493903E6DF27AA32791BE881276FE47A562A4FAC5335CC2BD21EBD488DBED137DFD288C87D4B56EED30B9A34AB295061EEEB0EE5E87112B615E010EA04DD29A3A0EE4FFD083E4A67DD320269D7EFE2AFB71E008279D28ECE96FC8274666925A0D3B42E58E4EFB621F3FDF1EF9987FD3A344FC496D0AFF92EE7216901559685E128B229A9D1561179DBAA0E08C086AB81120966875901295419E93FF5A73ABBCA65BBADB38AA627FE34CA63F8A0EE33DBDF7D2601FBD47A703786DF040D84EE16A3C78304EC38E4C9970129FF249353BE188CCC35F68D7BAB001A57734AC93CFBB85E48F6068AFA5F5C3897B3D219470283856416E1E256D526859DF5F440C6EAB7A86152429CD9719C132D6FD9926B3C69C55A0153B938ABCD31112C82A75BEF9A8B74B8316D61EF73D357B1F541B79B1A7E13FBDC019317A5FB76C8DC68BAFA3B8CCA73832178D01A298AFF65CABAAF18147507942EC8D9A15F2559A31872BC900D4685D2A6E279ED7B1220ED9DB5E3297CA4CA50179D93F07691B13B25C687942C1E2B50D78A4BD26D1912789247F1BAA82835852530E9A7CCAD49C1706C37A2E5262A1056C694AEB20D37AE7672051A6D1896D8E73C50F50F2A8675CFB6D35A7D68BE91E932CC51D85CA78560D135ABFB8EB36F980AE48826B932CC2AC2C8C1F3C1820ACEB3BB3E3084F19527D3A201C01683389E71ACC79AC5843AB2028B56897B90577BB31BDE84E6EBC26B88B151CC778A6B32EE9A2F6FE05842D632E709D409DD2B2D44FFDBCA91370A8E256920E71F8DF25B802766BEC7D614F035CA16045ED88E3FEC2D8DFB463F9FB0CBD7198F369306D352014777D2552651416FE35ACDA5622057CEC2787BAE8803ED784D71D661E2FEC67ED0963BC98FD5207C8640FCB132C63E89E648D01CDDBE942698A0B43E104D326608A021B0DD8F032FD915C34E0233CB673162B657D1FA00B25FEE1B2F14A3BB00E401A3CEAAD6F73D754CF4E1B6F890E82BD5C696A235ACF5FCFF26361B44151144DB231EDC51E46612AE8E4C6FA0C65C5113360E0F4C0E160A4960014D4785FE5ACCB1A4BFC20B966CD291F1E67B46CE04D4E41FC1AC2E13CABB8980114546825D2D4E7386CB7E6766911D23CE07A448921E7F6C79E3E7BA565D3977D46ED87C3A9FD3AB0C77ECBE8446819A498A146674B8670B1FFAFEBBD81AAFA6CDA9458129E3AF92D33EE0A591985828B3D1740C21FDE5E08DFCDD5CF0CFD5919EDF512FFAFC4E3EB85529DC38189600F3FA518710F0EDA7A0589FD72C77C7326F50C0F21995DA9862A7D2B9205B8701A0ED6E92E8057913AA9090433A08789912003BB950863C4CC9078978BD390C2B5DD3D54A3BB6F03CC3E2D8F218D0FD439DA10BB3524EA3948D095FFD3A8CA08AAE309C751BC2C1BB8C5C706C01AC1A9302CCD5AA9C43FA387AA7C23EF1E07E416E8C8670C81FFF314E554EBA6041D55DEB1B43D6A9180EE59CD68BE664AAA1EB13882D23FAF98191DFF594B661DBFE1CE59DE1AAE0448CE62A6E2848C05224ABBBFC78C7BEAB750DD012E16F3123B8BCE1889E1CFFA43829095774BC312C8C7704797531D020BE29E9B4A4637147E3C5B9A3A6D67B141B4CE0375BFC3E1A26B84F60100330600B10596843A4F17A861E4623C83A75C89259C1AFAE640D829CAAE9A0EE7D82E98503534C41155C12033F98510DE87086C0DBE69AD58DD635DAAFCDBB4C0AE4C915838AFEEF4F24367AD1B7D0973C30283ACD3E80BF236B56AAACB4DA8CA9CC812F62AEDF7E5EE1FE6A50D5AF849B8EAF90CDCD9623DE474B248EC1F3A3E3230EED1484A38CE390C9838D1FF542D7F34BA3A94073121D6913349F38A7BA4129A2620455D9EA4426C7B97A1550F14FB00066A5E05C7B7E8A6D5FAF7411FEB18EF65E85226FBA332EEA7148AB4076C2D53CD231EF6EE8FC5A79C36F8C8D1BE1AB4DFACE179A544AD4C8ABF375D797A82BC99414ED072A3B361DBADFE0E4E93D2E9EC8D0C21E4B7AB04D332608552D30474ED438E6A7F0DB05D4A649606DE526AE30FD5A1E76B909463852D9D4C1071AD6D1A1D5E1E7F5248D5A291E55A9C68E38F5D19138C874633D03B02A3C1BD4B46CF42F75884ECD7D7104F8894B22A80E5C3EBB8853818440F2604F810A17498DC11BEA29061EDF458A9EC1C5CAC28418758A11C3C0587B42F4ED2B4E43B9A1531F9FF2C02B8B2F65F49DD5D7EBEC992F2F6D78100FB74FFC6A58A9CE70136BF13127ECE08E3B732EAECEFA0868A26418B7E44ADE984D67FBC096DF8373D26DB165280F862AFCF8F51AD65722D911C8BC0155BF699418470423453EDACCCD53C586A916BE3C82A41D7350221680D6BD5F7D44F1DF59D2363902D427C0D4B45E0905AE48877B0D97E67B6004F0A9121914B8412B820D909BC25FDB7008B0A4853F16890E7D3E877056D37B356E44B0FF209E937D0F6A1D6C8568F659DE335328CC8C6C8B20C4525445E05966F06B92BEBA05CA68E7A0EF59F2B4F02EF2FEF7F5D07401CD0DE879597D12430F14E1BBA4E18EF55400085FCA175B4C02AADB6E5FE8E184439F68D7AC734DC7A97D68242C2068B1D34C617C98A2D8667CD34F8818494130582C57A4D97B75C552D6D2B29762BADABF9E775E1D55BE2FDA872F5CDE3C8EBC560B7DCA032DF15D56E300E5CDC823E8AEB3C35CA51A14A2F59A4A566AD1272BD0A766595721606282F29C7B06416B0AB096C4C591F9A2D495F3E3337D108C7AD2794F4051B41919249CDE0E0761F0CCCFF6BE5DD5FCA46C37A604B02E64F92D5AC2BC00BA6F1AD15C1FE1FF07FD6444947F3C944ED1200188C3228254EFA276A58D7F7165F494A89341015CA8D9F03F19BC6DFF099310009531E1ABE16F21C0F9C8CEE5491F8FEE37669D6953967C6889B8E02E0C3B8BF8BDBC755C9B0964F736AD2F5C2F5377324AB4656ECA8A8541C24F81BE146C72F717A9A841C7480C1A7BEDFD05D98576E121AE3C5C9C4AE092C688D75178170037ACADB2F44CA33E7975B63A096CC059361D4CBB5FED8501DFFBCC6B7F1ACEE4024A76109022A71B09DF6DB8EC31DDC84AF9120125A3CE044E514D28C653068CD4E6BBCE5A059A36263EFD7E70B56BC5D4D14142545062CC0FBB391EB8792F4AE0FB9B01CD7C73AB3CCE203FDCBF0D76C7AF2FFABC0B44184D7360D84CA9D29CB6459603809B09D73D009B898015F707E83D56F53C31F4F7CC1B160E874C2144432844911341B34BC16730D76F918B025308CA11A05389E2266E007777EA67A71A61471CAD0F7F0155C12BD01E1428280B0707664B2DCFFF2D782F3E82FE689FAFE91784B835C892BB28D0642B6824654E4B3A6B85D732B701C7939A75CE8E96D696E39F52AF214D1935DA31FC30E84290433101AD901EBF38FB6D59E6C992F517DBD91BA6E3BCFB01F7D04D7BBCE40A0A87363860FF616E4DCE34AB497D02199C5156BE5A44D4657B9143E1E11EE3DFD9E5526E4371AAED852F036EBD96F8B51BF87894017CDB0A4A706B2C5BF8F639D5CEC4706006B0DE3A1F10C39D953950D22821DCFCA96BB02D421F3B92CEA8815C4A7A6715918223DAB401936FE545EE94DE85B656B225532736DEC004E552696ECC8923E17A9A80B136C2B8A47890EE06FCB11DBAE067C93CADF37F3CB5BEDD0A0BCAEA0FCDF6868B6E83656D8C2DDAAC8C575630ED4F3456566951EE6DE25B487B6422EC2BA8EFB2738D6BF537B669DC132C8827FC3590CDD36C4B3ED0F1FEFF09C08191B1E553422560A502C21470050BEB5826165403B94D5F19B01B17723B75607403796B1E194E879D255BE6A34104D8AEBCD85AA23E7A644EE704C7C1436701A49364D04A88A6366B3206946E914DB711DEB99A764CC59A679F1D4DFA556925353C15DD0ACF91D66625944DF48F5071B3BA586803B61C2E5A01EA56683A88937A4C08A8CF57142A3C4A699CC07F489532761BE4CF2E7488DB1FC66CB84BA52A4CDCD4BD6187D947371DB2DCB11828F4ED76CC053DA3FC3E9CD50FB71970CE942881AC884F92BF9F23A18161FCD34E2F088752E93A1AFFC8D512B808287A0AF1691F7B1A7CD5C141172B2433FCE9B5EA44D73A5E5C2FA9C01F1FB3853CA6949D4171C8A073C0B8985475D41DD332A5FC476D9F1BBA2FA67D5604C3ED57246F53B0A778DE46AD8E83053A68B97BDF78581E2397C2FEB6E9CF241651C4E309E17D56F69F30530FA3A033E9391DDC2285AF27C438147B6241E34F4597D32411626E712909AB595234730B37A31FEC01FE0C21F5940EEE603BA081B7C01236393FD3B1B1B4C1690B0A1372BD1996F66EC65A23F33979438F70C9AD5BC51713FCC77CF4DE1304644860A70F7A44EEA171721BB681A9F5DE3B178C5F1B0EE934E28D6E0A4013C97DE45ECF41FE23D2FCE83E457A5ED12FC5DA034CC4615D06934D37F58257CDC9999F3AA3DA4AA45F8F61D5BD818788FEF8D04C26BCBFF07B865C000D7A56B8105F721CF12E2183FF0FC0857D5EEEEF0AB141A3089FBA9E9E4886B2C7FFDFC4D95A44FB3541527F7165F14E0B09DC9BF51254E06D157ED41E4D9CAADDE0D02F0A5A659939AF3140EC87D79872BB91ADBADF321C005E40B7AA96D9CF8C2E78546F04F590F648C1E93FF8092BC71CE26D6ACA4BC1293781B36AB7DBF5A65B133FDDA471D3C784E31A775349FAE7C0F4286D14AC942DDAE0AE894B940187F34D9C95FC014EA5920FE4D3C797D0E92D3187992A1493544139D87497FC3B08F7D86B7D60D66C4E6FAC5C88816A2EEF0B6724D6E46BE1743DF6AD564BCFD763F46271185195CF3847161DD0F806507F6E2673FDF2A3ED3DCD3FF60C4DD2320229EC396886D6653A39166C4C53A2D7E494855F3026C9536E95452C2DA77C5932A8991CE2B749DF5EA39A72FD3619013550E68D0378A666F03D36959C7A811328A3A266F415AD0529613DA43882BD0BC1D8EFCB566AFCBE32E0F0182653A15A3201DBC23BAA4947D033EA45E01FB77BAAF710F0A0417261A9DC1076FD8E5CC6D03FFDBA8229B978E89228409FC103BC9D87FF0351FD31C573B5663C9870132EA0555F233FF95F5C6FEDD9462A4245EF0F2578E294BF608EEC39BB275C192988C732776EFA6A240B63EEAB94D308D25BB2493B199F8E62868AF1493BF8513EC7F3C01F9A8ACE1F6D3187695DE3277A0B43957961D601B5DEC84647ADEA7FB37C1A009A8ECD29C745D2CEA2FF0839B544D5E9FB20541A7E54F9CD6735083EB029373CE44A911A818156EEB8C83F5C722E217E06E664A36DE2D7667A4C5E402AB487608075B851840C712EB6E281F2DF2F74C783FFA29301899BC7F8ABA0E99E1BF8825D5AAAE02180A79E43B96D40738ED2FA281250168151F9CF73EF2B56A2B3B33D0B7B62B439F603F254F6C4C96E1F96CB10224F18EAEF81FB08D870352375B9F94E6A9E060C282B475D617F96A4E9545676192538516279CDD8DCFE0558B1C2F1144D5E616D9DA9BEEE97A0A1A40000000000000000000000000000000000000000000000000000040712151F242D3100";
    verif_kats[0].PK = "75a8f4c956c0d7da6c7fe78fb03e722ed1fc4f2a5e2449600e616f61995a4a88babd92571c6802539c86367bac5d6c33ee7ad2f47331681daa2ecd3272a07c9888ef4fb3d7d7b5534d62d48db4e7aab9a3dcb6732cf5959d5acd4b258fd9aad057598db1a8503dd8f788f9b551423a93dec204c8a67890b533bdad3544e65dd2da8876e6803e5d77c6fa1f1c232ac0328c69650c63e23fd724496b95236b585f76fd7c949b0204ddf23e55c883c88b34a55b2d3b377de4122f9cbe78143efc7ab9d23b9867f5f939df336a025653b525d7f23586f82c3aad578883eddab3868a08115bd0c313ad31ff44f4f6b855025e5ff68b72c9d353ce54194914b266ef4d3f1f8740142a53d1c27bf5ef2d7e88402c565079247080ae0d07d6d7568fb887fe18bcfd8261ed2ef494c18a8e6b8a209781a4cd2cd32cf61ea4474e74aa20a22da5fd0b4955db1e2b9a6c3c38072c9042d2744a5810f3c3e9645b84dbfa7891f5bc4e41fddd2df1bacd84ae80bee0502cacac547fd6521aefcb4b95b58bcc194c6b5a4e5214018b6f2ba80f21122004ed559a86776826f3d777c25a283eada7bd2004b88e19d7b15fea24a153c08f0936e896ea2ed175c07a2cd40081d147087f8e7e8b56bd438f7dac54ba3a2d72556bacab5c6a6c8d632acf6e411e1e9299f2a2fd4c6519ac2262abe3874871039d177bffe6d167821f05e46393b1fcd5a2ce192183ff741b185280a379840c75b9ec706c1617db9224958572bef0158b000f6c5bce5066c4e311509efb92437c865ef4f6c2e8493a26ed8b2fd99adfc161a9059dff794ed52af6c83b7894fb2c79265468c230cddf36bfe6ebaf11463f0ef4ccc789ef23eecf3933638ac5ed3bfdc0122b791efd23d7c239bf969b886ec3626cf86b9d012c2809ea6ba63a4f8e77cbadb40f1a8b7c2b7ac21c00d3ac87d98e61ce6691a7f5b2351d80d8ed30b5a9006153a4878e517569f192f94f84bb9a4f35a45bb41ee126d93c19db43a981c57377dc9bce867a76f2c49d0d9e8801a1726c8eeb70f7ebdfac83e46a9cc2718502e590a9d70e82a9ccf56d33526c8e2575172c72e4259aa639999175827b93803c5b43e50c8833a80cc52a11b2c959b5572dea35924e12337bed0e92a4efda31e1e161b2b57b4828e9d95685e7db7ac795186a8b966f90caf876f405f1ee9d6459fbb2740783870fe6a5c3fe8036ed647bf544b88958c4f263409f56a61588d7d8bbb4073e7fd7c3c9e25006c97bc180435054414cefef80d77dd7dc81099f4bf565d4e891bd86368669faecd31f1f1a246c969838432715309aa45e8ed861517c13ac94602933a2cd3bfa06735e62c4beb652cb122579488ba8530bb5878787495cad696d7c5e1de65a66e4fbeeafaa259768ea2608ed25b5586ee1c06ceacd5510e4167f7aa4dbac15c68a2a71066096eb8f0fe6ae7345c2434a87d28bec35e506be01af27edf60752de9c9014b22de55778ac5010c780e79fcc357aa29326ec748bcc593e62e6dbc51ffb3f282033e8935d8ef7efff37ed6d1cdf5a204558773a1b8c7ecb87949013bdffd6e8e05c817e86dfb7b6298619870fe73e2b60992209207d94b856fd56f4c39ad937def57aeea0c832f54bf408755f3988a39ef871335bdc2169f675c95ea2658266e29e39fe97c0c2093e8a2eaa9db75a6a4fee8f6889be3a606c79956c24f3b560cce1c37161453868d9bbab0a87d85375126b6dc3e0d1f67b32a0006a8d3c705df2c6b03ba0fa2b9634c3b0869552a0dac3b21ecc8ba17b341c2210d0a23b5fd68bb1335ac96c3ef3701e0a2acd3890a4aebc908bc063bbf2ef3d50cf0f8da48f7ddeb86f9d773e544c70447041076e99c93db9d39780df774da35a0163da3ea50f17a69a214410736015a4abf71f43083324951fad485ebaf55de945f8c6efc3e8be26917e5a296050405a97fecbfd2625fc676ad1a9145bb8a9c1f1b3a46519f77da83c44d2861cad6a56ab01bf84f7709f0f5270ec550f6691c47e6b18f4b5b884118fd4af03d30460119322eaef583a15f00a561afc4985393ad53b681d41d469790a24bdc6056eb92dce833ab33581e08267cefbbc20676192a7608fb7e3422801d9351843b476263c0d1d5442613d6eb9924662b20bc213ca335a52a5f3cbcb8fca9d9164170c8928dd5d2eaf9290d82ea8ff7299e772de20567c79d6ebae9bf5834cad8d55acca5e9b22e9cd0942dd262f06d2b21c248838d8b76cac91e98fa4d5369fe26a609c2e6547c29137d45e4f4b08724df786511fbd75eb72dc72db2ff0b8d90461eead262feb1908f0605cf60b5f48733e3ee31b12eda1c220eecfca7160eae73da742aaa3408149ee255985ed681d733ab49771bbd77e344976ac45556a83cf5ea3a557d6f2d854af1396fe62bf2a582f3a252b9cbb00aff5e7a5daa0b44d3355374c70bc6117dbcf67cde2c025275a49105bf0d464b554761c8e0340fccfb2993728381f0a015dcc10d7a26970671ff41c6c12cff6e71e16a3763964042ab8ee7a1d9dd7dc8c73229061da4cf614d2f5336628ff9dc92a1a5fd33240ef00575d5008a2f1a632b7bb843ab18113b1f0975b6eca7abb6c18c2d17c9542b8ff6e99c186fcdaf6f0ab62dd37646277ad482d7f066c3c7678d5a9acc3c162c8ad3ea326ebcdd518240a6040b717dbe698f6e0e49f35741289a61f143bd0c2f33584733ea05c0f60321ace1874f0c2ff2730f729b9b20fcf64994719b95c0126af36e379afb8940ea28f69a43602a1009181547aa7f1c6b59bdfb5f010fba702e193d67af6a2d0277f474e504280eb8c565afe7696d8fed00cdd560536ea3959d2d7d1dbd702cd325ccde51cdf0c1af06b62089ceb523ab942a50a36e67c786b83f93c29b515cb56af23c5412c1b2ff1be9e01b53b6325c54f3e7fa5fb3f2d167bfe6f7aae10cd499486c74f26e76e8fc18e7fe42b09757222dddbaa0d97f88aa1f9fc0cf1c9f781b28abd0a7eb9334646829fddfc9f505ecd9bc8eddac160366bbc04aa2e62a7a209594a87f9e121dfe961da3adc7764dd63844b4fce43478d151fcda95ff1770b3d87a6727fc274d7ed11a1f0e286992e87dab4763cdc33027fb60d42a3065017214496e54c3d0ef5953254c02408d3ce807cdd58ffdce15af94762c4890f47f6215fbc28382f72c9346b4d74dd7c768a067ff6aa96e495dfa9d13470b6adc362bd8c442d77941438944521f67e85673c5ff373512909b8371dcde344cc8a602c33279033003c4b7bb51354b2e66c415e7cf3cd013004cc968be01a21d9104f92e9307d9d9581c2c125581739cf740dde7d530e22a3e08117559843a0edf0b6d576b4b528c8e21d00fe8814f357d63d0f4b091f4a9b4b3de3de2f3ddba9528f7c6e95433aea0ddc9077472572bc7f015542cbccac3db5ea7269cd97e060e3bfa854db263906946e6e5a973f355dd585da0d39603f52918804240f4c8a2640de27cf9cc53003201b6dc58a2ed125a52f46444938a93fecdfdbe504898fd127e70f9f1ae29eef61e6ac0d3b7c6a84561bff144eb78dfe9783f717be8381bf9458250424b61f095c1001be264376f4ba325ceff9bb4752cd3d8806870b5cfbfd252637364818ec11bff699cc10f3102fdd62a5b527ed7a";
    verif_kats[0].expected_RES = "89E8DA09EDD3600C15A06D5B5CBCA92CADF08F4313D0C0E2B23E24B329EEBD1D81DE6DEAE3F36797A494BA2121E0A274C3988770902E2CB325B79FD1C6ED2197";

    verif_kats[1].MSG = "ca393154ce0e065793750cbb96156c74eb704ed0f2ac97c1131f250f550e1efab980c2cb146960dd7c0b562a1f412c6b2cbd203e1f048c73376590bd39d7a969";
    verif_kats[1].SIG = "8A659F891085C42893C7523700527092698C1C191B0F187A493139A48BAF373B92B6E6D9D507A0BC0F9CA86226FE5589EA760E99F2D4E22378E4CA968A3E945F1D7F36F97F7C11CFA5CD67D63EFDFAE7DF68DCB8A3D6975673EBCED7D8ADBEE342F7B8E6F32E6420B520FD284F72DF044D322B15079150E6BC6FCBDD3EB6FB175238E3306069B4EB7EE239FFBAEDA41C704BC3F38280DFBC2EC22DC806357E4282F41D3C63FC9F6B3B0A02AA0BA960A45066424A59DE99D43934B48BBC28C8E30066214A1E13A967D5A5CFA25811C013D85BE5BD1490C44F2ED16D7594011AD2BBB4339914E650A604B907D8EAF80FF24A42B0DB618D53C14857344951A653170621A225A06F70D0329C3EA15798A28C1111C2E4902DE9C04C54525254792C5C0DF0668F2DE6F3D77CDA05605A7741A4BDAF5650A76E68BB8BE505CF1B4C18EB3C3820A7A90E69E5D170C87DF46C29F1E024987681A1D36D69ADC6879C0BF785A8139E2A857DD4A76B29963DD28ABFB9415D7010B54A496133E5BCEFBD9504C0A541A3AF30A97337B249F585F604580333D83FD453E109442E1E0E4E37105781F4FDB9590B05890538BB61414C3094E0E110116FBC25088F6E32131FFDF3E9AF8312D603E25B695D8F6D9918DB442BF60F2C4C8F395A7089208D4CC82A99AF093EE32C216BCCC4E799A0FC9A9BBA09FD372FDE10F0C448B4B9DB4631D03D9EBD8BFEF09D686DCA17D1B14459C0190C4CF9EB53F47F4E95768364CEB2A9A36CAB718BC483CBDDA9BF1AF881EA346EEF7BF245E09E08D3F355AFBB0B3F6420C725368E5DB7F6182CAB20C82D1363374FF9E18F444111923E94BCFCD236293F4E47C391184CE4EBCBE1716B1638B879F7D526A12C4990B552344570552E0647602D0BE13F4DFBC87C104D73760EC31EEB9C52AF2BE770D73CC4794A88B61F2619EA0AD19E90BA1BBA75F8892977F3935EB3273AE04038B94AE7C3932E10B4D45E24B5EA4E7F767ECB2E929CD0C48DD5BDEF58646A17A15961FE57E008DC1B5E5331C8D2E3CB3A3EBEDF405476D33A53D707A38E9CF5D9066B84DEB8AE8A75CD776877B5C44A90694A970614E7CA109BCA9B76DA126C402F814B8A2D22CE7C2F5CBDB70C8A0595F922341CF32307E5E69030072F91B32C29D1205F0D585ECD2862389A16ED461E0482F65B3063B093ECF46B603863FFC85800041650143D5871660DBA750F1102BAD4EFEB3DDEA86AC29D0510E00B5A811586102A667B76F997FD6F0A918782327CB374AAE591ABB6175AA15506141E54E622325DD65E4F4C8F69370C6D82F3BD06F80B04DFDEA8D547B1A2AFDE90DF654B37AED1F1DF080B24BAB6C3D337A25720AA73DC3E5CCA88F71078B5D3F2BA1812A593537171691DC313E21E9012ED9DECC6D20416F840E14712D6AFA552022C7B5EC578F42BAB2F77661B2C4754541252251B179FC765DD52A9556C650E795CB153B2BE5BC8AFA721F87BDD996F7A82BCE1955F163B6B951F837E5FFC758FA92AB83D472199DDC8942902713D15F5D1B57EED176AF6366FE11932507221963D8D332911407F04AB610DCF434688976EC347B2B6748515C82329A3A5D31BB3D5A73B0959184B1BA8799ECBBEC94B5B5DE2A794810AAC46D94E2210094ADE4807E9DA3F26327A32E019C52044D80CD2502E67FAAEF5087ABBAF93543BF9DC3D3544163C469952AF12670BB21CD946210E059DE868A52B34BE30BE951DC81092ECD0CC261803E25B7B56F963D58EC92399EC96E095721E2A4B1AE553C37C90CA8EEDB76FFD1CF7F0B7223E6BD68700D2B04626D12EFA1053C65BB14892C623C8872B006F8F654009AF571A6F91D83AC8E6A3260FF78F946A197035BB4AE04DDC9BF783D315EE35ACAD9BEA041E5C631D2C860D4402A865CD3D13E82A0158114B5F51D403A769277C0056C4C645B29177B79394B639074E85918E4D9244EE4C2FA2E1DA05903A516C5054B348FAAD38696DCA8214914241F658A0A659D36A96D96515D055C87B2E628F4FDE39E18C2D0F164DD1893F3E595F11B5463117BE1EB276328DB1073AE17EFF6419652840CF7F99B93703C1FDFD41102B02AA6BEDCFFBEABA28AA3BED6FA8EC790243679E629397E64384493598C433E5A34F1A96EDBB9697094D16F33F1344608E3122361B25EDB34AC763049F5EB9D21028553893659049AC318F6FB55B6FFB13D245F09A413D06C6D9ECE959C2FBA470EDB17A00B9432665A7AA223193075D7CA97B2298437F77F21775F8867270B9829CF8BD7CB76BE6C6E8F1036BDEE6E2DBED599836A43432876B44BE2930741CD934E5D0291A8457BF0A612B99D51D6CF4C412F5A156222AA1548AF136CCE6A57D3BD730D0B0A3410F4303187CC23E6032DDDEF14CC65B45671A8C0EE608881CDCD7F558ABEE9714F25D5C491068E3E278CA01209D96EB6EC8C679B21DA34AA9B494B4A67F2C742AEC06653FC66D4013557AD388E8EF21071FDF117102786D4F2DE16A68BD4380BD18558BB29FCE4FF761DC3D5DCF48289198B1DC586EFFF23FC9A89478217B37FB6F69CEB89EFF9DD0E045CDDC05A6582E277052E51C65C6DC5521E2F59B854694FA985D05E923D14BB7EF6AFE34E63F25DAB21F669AE6C6A9CC70BD8FD72D30C9224D6ADB2F5428193C6190BCF1C073B409B0C35B658ECA358C2B9D24D02E5F5926AD2329829926C3F39B0FD49BBA44A9D3C5966F07B4A06243AF5CA160DEB492E1EA4847FF4FD14CA75B40D125B48ABBFC3E5B764A19A1D491AF110D876FBA529D3B5D3A3E48686AA9AB26947F1FA93D9D40C3DBB36FF652C7A30A3ECC728E94583DFF9AF8A275886214B6AC055F3323B9AB25B3822DD0C2ED64B95E3DFD9E4F50D547BFC790694F38CFEC4146DBD8DFBAA2D78B2B3E11F340ADB8BEDDEDDCED867D584F67B9F3601A62F2660932901393486156B0D61FD6E6B459F5C01A485979797F1635687EF246C960D64C1A248145F5D1658C27D42F0169E71825EF9AD8893673A5D323A05D28E444660ABC4030BEF6C66EFCB057A9EA0684B1B64735728DE008A65E2FA43B84CE5FC39649AD06C92119DDA9C70DBA340FC4C27DACD809637D4FDB0634684C5936B009B5FC3FC7D9B09B29C70ECFF695D885A35C21EBFF236BCDBFED085F7B4E609626221571C8112F03748DD010FC97FADFCADCF825B0472254C026A0C5E83610E870F75988A7148F2BA399E5891164E59740BB41D6E6277C73B1412993F91C3E2DAB02A4F12C427ACAA14B21973C1D442C79D2F038AF9AC48A0D5E12EB82E234615BB8692DFEA8A98D83CA3DD9033D7C48B00A0731EB2DC01377184BE6F2D7DD697D44787C6A6053E6E628437FFA0419A0BEA50FBE52D6089A71B2E82D002EE1FBE6BB3108CE863A08E26890DBB769A417E8926950419D2A952E20AEA560EFD64A525B63E46D2604DBD2CA4EF862BD3096392D5455A21095CA663F886460F592BC75555FE9B13A00A8CFC9D6991488AC59CA87B8A33C472866F821D20F99BD228509F561458CEA2D7EC30048BB547E53DC48F1F976BBB304FBCD3F1DA708941A3B3EC3B7E9992ADF216FE127CD16E5E23B08A7E364704184F659DFBA2719E3C78CBE2F19CD4A84F12D5F60ACDB839DE814C52D30CB8B216A443B2F98225C4E18653CB36CFF848C0E07FD925570040E60B9810BBFA1FF2FC92A0F9EA3E3C74DC443D5363DBC576684182B13D573BEC531151F32F94C1CB54533ACCCDFE86DF79572044054713F3A83275D47B552CC7EEA9501DA6982CB81EDD982CDAE683C10EF122BAD67AA2B69E1BEA2F628880688ACC773ACC727B0B33B190EE05F3BF5523C610CAF7A838A7B9C3F185D44696649D354E1DB65D76832EE32BA1749716BC509AB60688164A030E06B5866968B3CD64E26950B0BC99517219AF04AF5B79EB593B0FE4EB497293A688741027F0725565677ACC6E9432901ECAFA14DD2611144AA5F4F0278DA0F9D7502ACCD271DEA06D6A89C42D473EBB50AB9087202E8ED9E4C1476B48445E3A7A3E022F32A220BF29B5442E41E0106D560EDB47BE768D620B13767EE72E0527D07270D2178608FCDF80284668CE9B74CF63DA78350CE9BC7CCF87B38FDD5C4EEA3CDA098282285D14B74072F07524B0E68EB7E780EC225D6EAECC1DB7610A757508D752E3AD82C5D838B72677FB78EC5D5C0A6010BFACC9AB90CD159280F440E886435FB8A525B8AF97469A8985211A83FEDBA6A06D713868D544F104994EE93EE0A3C42D5106B6765210583AB868BE1A5B9A0269757CAF882A4B3C2D4FCF8DC4F3BDD409684D17235763013D3939FB4BB9197175D6B25A966399FA0BD6486A63E4A20B91B987E955CDE99DED263A9EC0796BF3D14B2DFA3BEBCE7CED3E0953C02A44596B4623FB73F60C6BE64F0DECF9D555CEA95CE07C60AC56CC0C20D9E39AAD4B51D94682C0B09010E9BD1A8D24E1BBCE8FBDDD30980F03D67A6413B95C22EF21B4E889ED43F55D787E2CA0CE1B3E237B46BE54B65CCF93E05CB4D63141BFA54F90CCC5B239417A8AAD7A88FA7CCDE45B26D12A664F49A8154A3965FA8E3CAF276E35B6AF06D8F271CBC18C17253C0A7E21373E7CAE61F6088CDFA4FBB434B206D45A3B937DABC331342D39CEA1FB4C52FEBBA4F89136AEFEF338F021E4AA3E0E028539A5F126EA37A1456655311493CF992ECD7602E150A290EAD12C9041ABC57C13EFB1A3ADC7F3ADC7690C8217B85D2D9D92AF969EEE20960A74759FC0B91503A391A7CD57FFC822CCEB8CD555F27C463F486BA2AA96FB2776EB88714B3225C3690A108D14406D6BD6241EC15CCDDCE4FDEA4032A667641144716BE03D02B52BC002840882B9C377B2BE19CE16A49867CF236ADF14E3401DF348A642548D36E9FA1FE56CD02DDA2CC05A50E4BAB45174A8BBAF0DFD8A2662E96DCE4F823509B2FD9172C85C46F281EB9785D4C9810B7DDBDF984AAF2838D7C854CA47439D4D359A7CCFAD80D3BB18D843818A0F6476162AE74766C55F217E2F62230EF763A34B360C7AA6B3C531D6869800AA8D933B7BB0E63FC942DA2E9B194BC55FA64ADCA4DCA0A58E898C437CA9D1239F50D9CCC834D9DF1E6BCDF8EEA63609AFA46852324B31B96FE4A535083423D59560D1AFD42F3F3C57E98DB0629AAF087283DE6754276173D3BF388702E263022A30A224466433239E6F0FD13570C6B96C491151EF1916EDC7865E2ECDFA2CD5F32332E224757E27C6ECDCA51E34C498D42BF07C3A7A36B24EA3D0BE1D668BF5D011577068C05A8EF206660B3460B252B39F0BE21122CC46541C4F79148D6099F78B2F7D79A2C8E0477DC2D19E0DF277E2504ED60808553640BA21E2427D84CCEDACC2390901D4D263BFA2BFBE18596AD80DC44AF44E7B2D0F41FB9EA0890D718DE8F34201C1D018DD89616884291C14DCB0A3C985865DCEEEF58EB8593E1F7A7904E704653E74371F9C691BFA337A63C60CC1EC7F3FB0EB21BF8AD4E1029EFEFE5541A3447708D8268C70345620AFB46C5004D2C49996215EBC2D14302ECFEA6727A5D6BFD625FF858B8B0992F5B5DDADECD788777DCFFD17126BAF4109A74ED7A0E24E1F339DEF1E19C237D3CBBF070694E067C95FB08DF8C6F43B545DC4466C05E0B3748B3FF01742270F1CB619570E6EB8959E3E99D05A66BF2C37BEBE515AB6D3F495C397E636B9CBB9C111BF778508C73F190EA4CED77B8015E97F2F78EE087ED453ED48C6BE372452C22FADFA50A30BBF441FABF7D87698C6DE497F13723E3A5B6BE71783205AB2868CA3FA35AED4D3C73A0C34DD21972F693F0C47BA839F27FB406215DA997C65B4DDCE96C37EC416BCD378884831651D7CE60701B034C629D33C10B2F000134F1E84180AF6AD365B0AEC2D2E0A1B080DB26E9102CA17F82D7073523BA7CD0A8ADAA49ADD73F42A0B21CC6C70089AD15937F21B0935D77AF65BEA0CC5010874EB966BF29196100FFC274E359AD514ABF01B5FC21649B360BEF9B2A39034B9AE50DB4456B4C43DA6FDA72994A184D93C7134114BDA317B6AAC8F53D75D905F6EE49D6E7F5C48C6135B1BD9A88DA1FA35994EB775EAF760306B4915181BC51F61DF9361B6ED38FFFF4F0E66CB15EFDA30FF1DFA41AB8CC4515EBC7C2B47729261C1D08412D791354BB2431CC9296C2DDAF8982036E0B3A609651C53A2AA6E505CEA9AE27F02155EC21A0BF635BD63D9B145A655D48CF6E527698987FE67E76855D710DAA8BF19885DEE24448B8AEECF685FA241ECFCFEE3CF75E54E762085AC0228FBB8C87A2ACB57B3DFD585E8C8CDCD8EC03E34C290A521EBA4CE37B9E1F446B9F4A1B70666DC9705D6ADD69FC206B817BB73A87F4DAC204D1151E24B8FCF7F6EA0DD84D57B85FCFBDFAFF66C0CA32A0251D5CDF19252B2D685BBD746DD2A5E8263B5154838586B5CFD146587BB3CDD9F30F141B38575E95A7EC9EC0E4E6F412475863B9DCE3375B6677828690FB6699C1CC0C4D8290B5BCC0F500000000000000000000000000000000000A111A1F262E323A00";
    verif_kats[1].PK = "D7B1AE0B7AC9DEBF3236824CA48B49A5FF417C11FE65C667716FBAA44D3DD620F5EBDF9D49AF3B711F815E9BB80488C8F3106EC723E7CEE24F1408D73787A54AD9185B8A7E331F6085371C71C5A94A64B11AB9C2C05D1AB0AB8E2F6DE7A10E3562C28D10C563C57517688ECFCD7D2C5103511CEEB38C17DB88D256DFB1282A2A8D668543C2A5D44E01419F2FE79A9CF7708EEBADAE74956B0715E9FEC122CD98163DE1B961A79C343655957EB046E13CDF26C3E24D625F751D28E8B08BAAAAA2FD10D8071CFE63C875E129B290B2FD263D306D502AEDF01423A182DC1608B392283D0C5A11EA510048EC026E3D53A8F6124BA59929C7DB8AD898A6277218738C1FA2E51B338E7F2B7BBC45F5AB90A911C62608B663FD5DBD157BDF4C62CDDC3A82D8C07D70C896B37B56CC307905BE965B17EE996A1420044941F3FFBDCC6398E3AC716C78DC558DB07EC6AB6B2BAE75F2C8EE5A27BA0109E1993017D98B42933D19D9E0DE56D743E6CC681E2179A6972DB9EDC51902E6527A3A9D7C53B66AF3BA37D62684C0CE046798EC4CCE74224A1161E8F61AD01D44814E34ED69A77413414CCD597588964CD1D9824E50BB818928CDCE1FA35D470101EFD1664AB86A4C1FFCB2E51CDF2072BD8BDFBA7440BD9CB8643D5D8B1833B1771FF48DC532BE02D57181CBF38BCAAC0302E0B499DB4176B967973201E21B6E0E4D5ACCB65F1DF56E3D855F7AD2DB23CD0F838DAC241455A085BFE125FFB2526C3A71DB0EA64E756E0A5BCEB7992B10518AD366DBA6031AE43F4AC033129BA2A206ED17FECCA6747E5F350E0791DD0656125E682CFF2C0176F6A6BADFDAAEA474702BB1A60B4169F506977C693CB34DBA3010A0D26A5E6C287907E5CA1714A93890D9913D86EBC5900682CFAA0CF01573369AF40708F3CC83DF996CA12530B54958A288F58CF0D95C61D5E689ED2208E4A1AE20828D1098F894578E2C6FD1841A583954B037B7DB54DAFB11E6D8F38A7A091D777B36A29F90744C11D4DE7DFDD37E9E494E73C2920DCA5D8A377DA84148F0836C88D472FFD371402DE5A990D3E374F9478B834FCA975D261E79F9024DCD70DBDA745C776678C17B62353CD93A6380B849BE5680B679ACB0113C004A616D8E3208F89A52264319F973BA345E16AA40825D14D30FB179E8EDAF525AF8BAF56FBD44C97E0A3191C4D9A3DB9D4F9291BEC065988D82D39A5284F435CC2BBFE76367AC78E9768A12AC88F268157ACEFCC0FEA6BEF6E520A3603AFC090DC7D922D779B805AA38FB31FD95D656EF5DF3620122CA83DF5E83051CBCC2E6767A9005DF0D65DCD0863A3B6DDAA9357BF31D9E370A027458E687F6FB159935101ED576CC1A1965B51F1B46856C070F3EECA68D55DE610111BD831D34CAB4BBA7CBEA57065E27C2E2A075D2F301BF6B795CDD8C91A8610DC72E495A90419E58BACDAB419DE6CA5A06498E6EA382EC2CC284DEBF0AC7D52417CA1310484EE64C0C8385839D66A48821BC099BE9C267E0BDEBAAEDF2FED4C8D5C8FA38ADBD77B153991516C444B5D9F7FB01EA442B3F603F7285896C612B9332DDBA545B8342D9E553E7AB2C88A320F9206F9C72FE3CBFA15EC12541EED585484D9E7E0A97B44BFBFB66C48518BC31543C680A7D320424BB0A22697FE255E4787498F998812C712CF20DBE71750472C51D4AC501ABDDE8B90CA21476383E861721554A9E667360E030B02563E51973AE326BD3F8B9BED05272845B9CAED94188989624D70FFE5C6758A6BF6E225C641A3B71AED6F2844778C4BA844940544D8C8AB1D6556737E995EC517F66A60B616BA243E1739CB63443011A91E704210637807B72A993EECCB0C9719CD2FD3480FE45A4B329E7FDF51CC8FE9D136381A2DA3691AAABC604AF98465EF36FAB8C2C71CB9BD1C6D48BFFB072206903C6A41516212ABDD40206583ED0F66AED210023B19DAD522ADFE6E31586188566B7C64FDA5BC850691C75112FD5392CB18E5B1C2A0BC79A5FA757C5463F134980F2A203A93F759F3FD3AC4A17C71C5C6E428AB13DA82F3A52F45FEF60C7277EE256424542309C371B33CA9D1865E9F52D839FA9E578187B6D0C7390DB1715596ED24250AEB7968BBC9C5B77A73BC9B2C777E49B73F918D13BACF546942FF5070B760C1E624DB603DE558787F6BDB326B3C93165AEBE0B818A943FEB8B2DD72D8180917B739789B533FE057D3154159B0ABD67B60FF681E011E152BE6749F296E778461277F5AFE8BDF28AC56DAC78745545E3C20C8639BB76AAA76500E799078E59650FC82A0CB2B28A05DBF574CD9A50AB041D494A389D4DD779814A2B24ADF580880E95BC21DCCA392CA6CF7E9A50A3D80B5E6855A0426182489090BB82F1EA2150016B4B3EDD9FA3A2F8D85AD61AC2807BD814E5462545B82388A2CD33F310E316D4815F8812AC924FABDABE7E696E0FAFF17546F359430461053031D31BF20FBEF05A6EDFE9720E9BF2DCFE15D83A597B3BDC52714778176C3823364B383B61F5ADEEB770C3D1FE161407D697B6201D5F5B1121D034A6157E46F81342ABEE5D7BBB8977F6209219BA4B8DE936EC87054132CAC3FC65666199F48C20E2FD56B08D04CCD4CFECECE2BD1C65ADC9D0B8F26E5DD582845B761350A3A8E6179105B7906EA2DF4CC3C21402F0FD5ED1854A11CB59262819DF514CEC51C026A2AB9481AB229FE42B3A0494FCEC6C2F6AC160742254DAE4E4CEB4BCBD288108A71805EE27B994BC919BBCBFAE1E3436EBD6AAC2A56ACC37DA6D39B52266FD3A6B1331BFE9BDEDE19B6227575662CBD6DDC5049E205F30272C151BC0CC00E3A2EC4A0E012FCDDE6C51FC33A18C297F86AE61803B21346040099BE7B5F1527E9D648426F1A06D8F8F74DB968D439C04660B8B14EA5BFF205E273283FB1B40B47012E718C50C7E899533E591B54F8D0631181962EF810298B0C29414882E51B073B19BF1C49A893E6B541D61AA48E2EC909102C954FF63E81C40B61BEA01D642B869002D6D8BB1DD28090DB3CBCF1AF7FD0A17108C3842C12B4B55B741C28E303863F74B6A1998D18A7952CA6F1A6F83751A5550EB32A0F9218ACF9945CCB1181AEC15D750B74E6A6B170A6DFBFC7A09EA13089B6906CDDD285835D841C2F27F380FDA69A0679FF94715861146C9EA97A728E1FC7A7AC23FFCF8150F94DBD64F47BE44207903C64F2645DC7D4963CA94D0B97E395341C8EE2D52D015446F972415A5B651289274F57D55705B8152ED2948F8BFC84D7DBB127F30ACF4AE91C05C8D5C964992A4E6E8DE6B569F4E36C5B846A85544916DBBDFF6C9250C91B9523D5EDAC17505D6BEBBBC8111E89AB795298CBA5A0E25450EB73DCDEB643C051133408DA8F3D6B47C1AE23F1B010473AD0A2F62E63D05800BF9FB05DDB1040268A0D4F0EEA7AD172EF547A9685C4BA4AC0D719E607E96D4D20314153A366029A81AB826BD5235228AA2230C6C0DE15232F7DF8330536A5A156801ACC2F20BAD0DA972A9FB2B4566B48F648A9F870DE8181484DFE57530A8EB0E5C214C418224699824CAE98FBAFFADC7C9DDAF635ACB7C92B2113480FC110E1D43B6DDE1A755C4E11F197E7C8CFA38195774B65DB88FE7EFE0839C22617E0FE33139EFCE9342D2CE72616CDD58D0316C1694";
    verif_kats[1].expected_RES = "8A659F891085C42893C7523700527092698C1C191B0F187A493139A48BAF373B92B6E6D9D507A0BC0F9CA86226FE5589EA760E99F2D4E22378E4CA968A3E945F";
    
    verif_kats[2].MSG = "9433ddf6e491cbf5cb03720b542e432f868bc7b5a0bbafd914f210c3a9d145953c6532b8212660ff219cb0bd283c6c25501aee58ef4201916e7671f92b759f21";
    verif_kats[2].SIG = "9C5EFBD8FC4BC59259C5528538F9546FC47C6ADA017628AD039E841F3EEB41078CFEAFE6BCA288F8A1DBC40A0A8DD61D7CA0C5DCD435267B4352CA2E2F3BD346CC790FE55DF82A25C3F23D2D64B4A8970C1277A2522744027C90F0FA18BF22E49C1AE5E589129337505AB9ED4318F756911ECAB97C5E0343EAD34BA7B6B89DCC130903E9E0902941B58213C94C19CCB36033D514A628B3E99D819452A9298A76DF24407CCB332C55FAEC61CAB4C99D63586DEEF80323B8DC05EE160177046D298EBE7C7E07EE5570F6E4C95EA9F5FA6A72EE55FA7ADDBB09BFC096F6D544BEDD75DD1702203396E149C846D66B846CEA8A7718A627122ED3DA6E25A47887958A97A28F5A84A7B9E608A0D929CC0B48329ED824B2B39EAE56F20192F9BAC700C2DADB42BAD7210A76034CAB87576698AD61FC4FDE9A29193ECF2BD6FA5741143FF6D5DA8C125FA336BDB627C8ECFB327065C027408561685836107CFC2DD755E7933A2560B8CA5A13A5972C0F3CD1FABE9D1D31ED52E63EAB7C6F30D49911EE8435E1D58F42D24983484F62C6324CCA3AEF6279752CC429657C80E59D2CA789D82070CA167143B407290B373D5AE0F32715DA5040FDB844BB8B1B388E5131D5ED474004FCB10EEFA799CDD494397EB43DA9B69CE5468C13DB7E70E56A974B8EBB8636E62301161EE9CD92A61B9C00C389C784DC48EB29C3E3C03C13FDD841B6D5776583FFF2E143BA8279ACABD9B33B598CAED53EEF93333AD2076C5D4AC55625EE6888D67838B3FAE33068EE735F65BFFB8ED36A75071143D0DCDAECB0EA4BC1997778A6E919847B2127EFC49860DF42DB656681B115E7CA402D7395A3356957C9F63F6B53D7DD9AD681AFAD26A95B3844B042966B29961F2CAD3AE1B392C0F6E444F5F28F9D80302BE5AF3A450FF674ADEA63B72EA1D5E7C864BAAF1B1B2F6C65DC25073073AFBDE65BBD82C4EDFDA5FAB7C5639A5E79F4CA17143C4767A13AC4CD1942A1FDCE95F832577457FDEDA9FA8BD6CD91BEC05EA2AF3E77DDA26C233341147513E2E1E66079F6FBEDFB82B9C426516DE1AB27BC99C52EA86D16311AB303489693BAE687CA4FAF7FE5FF3E66D1B4509947C6A3AC8D2706C016BE4A75C64D0CB9F619B0E9310052D3A7DAA467698F54C043123316FB07CB095D389FAA0D643D9C68BEBDA18D3F26BDCF50C58271297F556C5F69E0F900C47E40BD22B9EC8F5762BDA9B6351817A93523B8C5AC863B8CA50E16798578F19DD85C80DD97ECF158944ED3874EAE1E4401B44FDB28053E4458B06B6A51C44635414CE5255C038FDD00B1777A12D52738298647E10B2C24A56932676305370B7FF2290D3907E1501CE17B67149CC83C19DC90BE28CD2BAFBB6FF08293FC2F0CA70B9083517F5BEA55BAC22BF1ABBB940E522916ADDACCF9B0BC1B2ADA06B3399F5908B6B517454FD84207A83C0813F1AC6802096DED339A162892FD2DA66B64C0E756360EA2A6D0DB794D5EBD44AE81263229F78F90543172758228F563CAE50C02B0E8918871D6F213A262B5C44D0EA31CABC478770B408A91FC7DB8E4A842E1C631951263BF836A338DA967582F4086D4A3BF47EDC57DBD6879D675322548705462912173BC8278FCAD7B546F9B9F73852724382A29F3904A06C8BC2E24BC0C6D3897A811A78EDEED0B8F8DEEE869542F936C7FF3AC0D67E55C95AB1C7A5F23AA1B989FCF97CCD2AE097A6E8548D97B0A76CBB2DFCCAB0C7D1AC9EBD3A8EB8F411A5712DCEFC79E9CFD3D69AF856E93925239FC666C7FF02518BABC50E8298766E953F95C2557637546DC7FA1B80E994F4EF93336122BBE707CEE4B7C2E875D2D1E14065A8636645A374D543E42586E4BBBA52D94E3EC1687C0488379A53C8DB5F409630586319033A06F7B21E382148906D16144FF8990B94FD90D4E85A729302410B89F121258033A7DA98883B50DB5E89CC9655CDFF8E9F041A075B7C742BEA13E36A83C5CDE0120BE9C59D50A0496A862432A82FC645D33C174DE11510873FE541DEA335E8054A0B193574CDE4E20CAB6E7731A1A28DED03844B3C76B9362565B332140F91AE84016758A0C4AA7ED931A509047A5F1F2E71DACC724808E8B30C96C5C1984FF406B3667937E7E9DA309B6A374DEE6E2C91CF7FD8F4459D4AE9D6C27310EDBB99390F897CC98D5A2051E848E8DD0BCCCC382FDB2DC8E4A4C1B5E6A582DA10C31B219E9670CFC53BB36EBCA29C6DF49E42B1AA34644FF5AA6C290EAC68938236913B8A8F970AF0A9A4FE56B2B441026ADAAA67E1BDB81D9FF9761D76E44CA7AC39B127048EBEDD8A2D41ACD9F559F2D0F575DBA0CAB52F8FE5E6031625DDEA9F363EE4CAEA36F4B6FB71CD079039867D22D089F4502A53B718A504F5CE1D0D16BDCA8860CD20D4F55A3D29EA7F7DB73AED014861A8C8E41EB39E3DAC98757EE6C3235673DEF318675D9E686FE85DEF0A3F38689751195460FF9BC8357191FB7CEB7A3F17C2FB1716301C5AA9550209CF8EFEF4A54E92FB41B1F962751EFE7A0C94B387F1DCD09DFFB76DCBE9B10D9436157C7B6755BD34321C99AB84335792EEC3730ACBD54E88AE9C0BF78072DF12ECD51175D4EC80EA45B2723BA6B9D4F5F7786A6F278078BC9D0FE09B4144FDFAEB86ED68A67609CE4CF3CE14B83D984007DA1986CB8488C0981C1D796B874DD70810601328E3CB1A72AFAC867022CDF07469CDFC1014899FE9BCE106FAFE9F909D4A25A886CF7EBCE107F52B2048A5D0A6ECA24532CBFAB0712B92EF7A2CB50EB15B2F9FD3FB0541A25E2DE4198202E9DB4B36012B2035F4F0FBC15CC6F121ACC19359A49381FDBCF74F46D80661996DBBE0D530B369BE69E0CA180D3CB9543AB8E7BA2C7BAB67C7B02DDA2BC9D070A60655A9FB0F90E6468F7502EFE170871FC0E27D43C3945A292BCF9BC01A3FDDEFD87E4BA46D915D918622998EAF3F64C3434E39B201921811D67F99F964DA3A831D6407F1C8C5311557E6D9FB83D55A03F19E6ADB056A1E965D90D1AD03F9B8588DBDD78FCEF81DC190944AD7FF4B9D1ADCBA06666649E5D8276D513FB7E148F3EBD555E0361A9D204202BE359BF4E5FB7A088C472EB0268323CADC8D5CF4E74BD9DADEF65A0395C26D57CCAD179257BBAA1C4D39B755CD3552C2A5A0C53ABC114AF180781F11AC83E7A5FCF7FD5A977A6223F6D779D2982B1E82CD6936CE4E29A6C5BF88D474F6FB163C6BF54F8C19FD556E368E71776048FDB3BF51E54FA2814DEDDA42FFC48A00516CF304CD8C6171922BAECDCC8779B43B73D8BA39E3C04C22745C61B7D92EEB8BF28C202375BF9B8801408F036685D0F04A11E50969BD235412443C4503560922750CB2BE179E4C9BDA51FC290ECBB5F51BA7CD060F6EDD70CCAC48AAE5E05E070A01874605CFAA6A5844B3C20AB989F6AA03DC0E9C5D046EBE0A819DD770849BB0039A1600AB455F46A0A6E11FBFF35CC06B4A87099B07F7C62997F0FC4BBD46F9A0001F031B58D2C1AC8C1B91ACD3BA2E3970B1AF0D11DB275C898A7A340BF0820F81370E957590F0E513A0D128325BE86C84BC61815BA37136BAEE6F94E0D0350758DF89B25CEC22D36515723C90B697333359AC830D4CA418859A42255163761642B84704DFA6E0C835560BDCE67E1D5424876053BF05B7B8310E0BB46299F3CCD677F8C67596FA268368463870DDD7F06347E8BB28BC7E3EA10ED6BF20A6939225DAEA03BF52D957990EB0A8DFCF403E67D1EA6EE6C48CAD03580883D0086546A8ABA936BD6C837E07EBD971245FAD5213EB5CC73AC6632051F5CBD5FC35F143BD8A30E4CCE9CCD9514626B986F2AA0787CDB0CF797623C41C6786A4D8F39C6749EFC1F06E968692C8B67ED4032200DA35A1C2CF393CF1851A184891F15EBA55560D12EDE777CBF5F95AAA638BE56977A0611E004C82ADB6F95906A3949BDC01683988348D3F5A47BC0BBCE22F7F147C429EB8B9E2FEB013AB6D20562B3E2856D4767AF8F8DEA16FC75815D9D25AC13795BF976E41FF3EC1599F36BD913E7E2D9AB5ABE7FB6FCF2CBA652CA00C3D84DB05C4BCCE42735822825E3DB5580075CEDA00F0F06500413EE11733C8C1B7B14680FA368EED79F118BE06E8373168B83821A2EE66349473CB0C36B16C4A00EBF9247B9E187E8CB4CC2429F3509D91875CEF69AA95552299EC7EB7947D6F1AA41A87B8DFD40F4F3D2465D7D1B26F0C4568448897115C4C3D007EB35270AA60CF47740F193A920291ED247FE5C67780F510FDC23A16DB4D1F56E4DA799EF2245BC2EBACC2D6B5564758F33A81E1BEB3075235AA6B132BDB0EECC4F98604138700D3D36C5B952F84CB50820805E8DD2D46E7ECE54B2EEE4025E158743C0D9422715ABDB76934237BD743ADA2795F5881B1A4139A371156C05830BB656A0D5571B419894D52CAD68E03C64CC33EE70F90819CE89A91CCA0F5ACF1594659DD195C8140E02D0249EE10BAF3C8068B765188627DAC302ABFC5A0B30AAD53F476C8E8A201CB5FBF85055D727894EFB3EF70C991A2D9D6C411923E456F4F8417705F042E890AD69AEFBE5E9EF5C0307FB1A99CE9E99C7830A383AD703503D5D847D703150920C423BC0A2CAE2A8E16F1FF30C932240F5B9239A4A3D4E56AFCCDC3A06E74FD5930B336052F9BB6029AAF9C9718AC62FF8352088CC6833D5F97352B4176463D58CE514D458CC5EE2B99E84CDB24F760EF7C737FA0F762FF4544BFAC078D4494C0BE2769EBB872802590E21E94599257E9452161968B6C2F8FCCB8241A861CBED00D2C38C3438A8A5BBC44C533B9B8BBF6E4F9DF7180BEF52062A465BA266B97021D16BF0FF8E29044F1D13798F47FA12791232E969484F729C699F7DDEFBE97E5ACA8FB900943E2EF04CEF3923DB07B9AD1D2880656BFBB365CFF326834F651A9A72181AE1AF6D9DC7FDBDE84F7D271984F948B8B963567F548E6E00C1648EFA7514E072C603450FACDA79B6827ECCDF9E607E9B2229F4976D5E7A3F3E1415854F2BE29A585B23FEAB97EF227BADC65206F8325FCC362A00AAD7B8187B61BE1AD29970EED3D6434D34AA81D6AFD4AAEA7CC5E74B43433FACE7E078ED44F84008D7CA3BFC44DCFD87E27F728FC2C7CCED887DC03D875305E266FFD83CDC31FBD75D17D94192BF7CE72259C37F83B2F47AD244A77E26B07B014A5F45003A433E1703E850D6BF96129079BDC684EB34081E43BB2020A52FBCEC34C9F035DCA3A66B152849D34B8E5BD492E06FB3F96145C52C56413F68101E609C93DD58362D24F4C849DB5209487FB47CC05A104C6E55E4F275A66ADFF772C84BD9B5651789982205367085DF95EE12B8CCC0CC6E442F98215A5C37952A732DA0E779333E1D35F75DA0F56162400BE8ECDC67F554AFF2A791C7B67859F1BC913F934A62CBFEC106841AAE74E88737E9C2C26305A32F5D7289BF25787C3C43909C175F40B895F3D8E34BACAC56F6406AF5F3F1AC28707099F68D72C841417AFE98F6450A46FDF89DA5909A3F1AD6CD16D6530396D991B6502D137A13BD91ED9A9461BDAA264746619FB4FA93B843580C68AAF80AED82577D16CC4E354F9D90EFE35F0A45ACA7D39831443448091B7308164D49255BC12FAA901E7BB0B98664C58B5DEE3820BC3497F0086B8346885403502886329442C71E51F7BC2759DB3E93F2193F74B5D923C5278D1CB41B6943E7F09FC36937A7E9DFEE6D5F20AA67C416123B66E7BA8E370DBC11755F912B65D16E29E4F3EC01ABAB2CC40BEF9286C7565806815824C3A4BA8BB3430D4DAE5EA46EEFFDE0BEC592EB00776E06D29D76A7A8ED633429574C9F9515C149181B9BE8489840B486C29213964FD8058497424832A4D221964C344AD9731849B654D395C18F2117CC3DF86B8BB37CA65BE7504A3FC27C9EA0EA49893BEA01028751C51826163AA95224ED6FD7152FB0ACB25C38017EA5FB6267CEF654BDABC122319D439B6173DE4538DC5118269CFFDD446351E74811FDEB87D3632C4D2EEF56AC06AD5B6C339F15BCC6898E36DDAF4B6A5ED83C37ED5C0B9E67372C1422302F9089452EEF0AE1D53A81200A44C6856ACADB838015B18932E682A6F7B2FA6CC9943F63469AFC460DAF780A472F31ED748AEB194CDEC5768B1B343AE64AD65985F84B5FDB0C98BB231B86D99DDD9C1668AE4F333450A713AA35FD96614EBA5EB3400681653327698445866C05347C84AC8A265930D486F08727633CE13FA0C844D3821F5727FBB3200AFCD51302E199B80F4447868E425961B19C8D649057B4FEFCF10EFB016670503848A1909868460E6429C6DC725E2FB5A73006F929D8F71DEA23B527AAAD638180E4339E82C9AADA5D06B8ADD5BFB077184FA270854B613A639084E6CBFC6253011D07F8F045CC391DB45CAE21DA014B3D67B9F55E6B04212243577086949CB71C1D7A818B8DBCE818254E7E85899BB1133235518B97D4DFEBEC036BACCDE0F6FD010F687F929EBBCCD7DBDFEB03579397A0C3C4D1E60B103D8EB7EA00000000000A121A242B37404600";
    verif_kats[2].PK = "58E3563D36F5D0492030B6E5AA317FD727165ED2F494FF5EE45F7E395045C87E4B5709DFA6E7688B11B81F70BA940DFE52729C62AC9C8D56B0A93D2D2EBF4347144EFBFCAE4BF801CFB1BB6570A8A58C27602F44DE8399E1EF6281B84DB2614F4DE383BCF4573F411FF97CA729BD3503FB2F91F5F778581E89A8A44E3C3C3A86893E78F991B7A7FDADBA06C938A8FFB66F58CE9B584FC5DA89190BA94E896784834914A4240BD8143E1A12BB78036168B09D1E4BD274FEB8084EAF2913617D2A1C6BE16B54224C552B7D410A831941EB25AB9ADEF774A1F73FCF1436D428E051C23B2C7B08CA788B5A70768FE2B6B202139177A153867A236A9FC9CEA37F47FB7E2FF30972DE89C0850DD7B38AC0F855BBE607FDCEC0E4A32E7928450EB1A571357AB0E137830379F9BC7AB2D8D25C3C59E56229A4DFB1B28BD9B7D8A0B5FFECFBADF3D24EE4E15CBF34D6E771AEE04CB3EF866083FAE94A7BA0853AF896B1438FFA79079DBA05ED1326479B79EF1B770057907CE068B3A62170936F42DEA21E596710A0975BEBB86D605A8A1A4612E47F9E60678602080C57D07451D6F207DAC1D55444892DFC4783FD0ED05DC61054D1E5E234D11AE559C35EAA3A5F6F2EAC9F908600FF2229F188B3C7C3488C88C891A0016198F6DDC951DEC5BA79D217A7779D18938536B8A049A8E418E1A73B77490A8A11A7FC28F100D3F706EB490AC59E38D39F30BF632B458F4CEF494D5132D6C74864737D05AB0AC85C34C91A19E4BC065EFE5BB4F27718D9FFA0431E5619F447CB8C92111EA5AD8104C57C47E5BA02985D0DFDEB9BC9A6FACAAF57F4BE0BA680BF83308306BA43838F7EB9A8ED5F1384134902DE002705100E6785B2DA943ED591CAD0A085A850838E10AE9889FFC1CD2941E1899E1A26CA56CB7480D260B217798056D35EA62BD55F159CF0FC363A4F325235ACC231BCAE18E89EB70A6970B2EC08DB004961FE951F8ED294D7D68CA6DB402325D054A47D17FF5B38734298B99278273021F165817E7805D581A0B9E40D507CC89D543F7A1B718820B1F8414AD6946B1AF7BC3AC1A520312240C0B499CF6B2742508356F9C366980BB1894D343E1BB24F06EB81CCCF5CAD59158FFD2C0D5E0019A839EF8AAF32292C33E32F6454BC03F7CE05D157BD875210A4276EE7C828291BD5AD5D545AE4711FF0C1332AFC7D716D104344E88BE87124ABD94216405A370AD8097D80879DDE60CB1F70B8F2230CD81D719EBF1C5C1D6EE965A85CB8C9982CF1625BC69B0C89D5D4207AD037DB73A929F024DDCC2306CAFBA0FF819CA596EA988A366901172C153D7D2A467FA1AC7E738F3335C1A2008181A8EF3064227FE7E72DACF26BB28816BBECFB8224167224BD37C5B55BCBA256C9CBE8B18FF4C36EE6A1EF091A714416E91DB1D638592D0FAD1DA51085D36D12B1255884B849B2B6C661A9FACBBBD67EEE7BF27CEF998FEC1CBA2E5EBD5361B429D509EBFC6CB2DDEC67B6DC69884A342D4A6C6D8001E9652A1486B5360A17BBF3A47DE94D1A32A5E2602FAF1A41B5908F67E9832382E87C9D432A3B8B6E230A58EA733F980488491E7043F327160FCB6D34383FEE41FE7DB76D5BA72B3DF23034E648E8ADAF8D53E1F63403A62CAF6AB88CDBDDEC39E9AA4233E3D335DC890DB9454CDFDED997B292562B5B001451729C833627E9FAC08097FDBB64464CE6B4C0D33FE64987373951F2E3E19E7CE119A82C2529C244BA56C7BA3C703CD7C940759403829A505A635B4401AAC9A8A9C76EB375F6069D6C3FB6511E20F1E9F1B40EC3CD47CB90B638329F17E1A3D9CC45769AE2E6CFD9284C11F4B0892BEA676F9B09CAA8E83CE7B7648546FBA7E7A8B9580ECCEA43FE330A0F1520F5933164F524CA22EBA3889A51D184885E515CEF8B35E65DB4DFD90D8D4FA1FBD0F7F0936E55643905AC144175A27F189865C011D8570E2A57392A521C6C38DD7CE0D3FB5FB4C34FDA41645E5BB32DF8100507B8C0B33846D12C5878D5AA05B86E4D83718B5158E67B4D8CEAFEAAD3760599C63A0594B64E21DE4C1734AFC875005B798550F02D1203D94202AF189F140D3729733C276DBD47DBCC0B427CC113A38382E4044B74333D6EFE559FA327F9EB5DA8CFAA99B882EE97280E7A909E4B23A0D35CA8164440B71699D82623BD542ACF364C6D74E4D8D79A0C293629474B5D8A05D3408423A17B9045E9A3A6245D4F123DA541FB8FC8C5BFDC3E6BC508B823DB3EA81D1529558416E720346DEC470E5A7FDF7720893EC139DF5B8A7664ABA3FDE76AEEC0EED445850B5FE0F81FB3D0CB9BFC1432EF66FB8960E4601B50FCF176AAB7AE4C0E9328CBD5ADB4D8DD89DB72B0221382D96C04A8F511659D62FB268D781EB68962D2167806C73916CD66DF16E9CB7A1C25C794953FC3C87326AC3195E6285FE5076C35A56F24E7583E985D51F8EE8CF24AB0E78F2873E426C20B94D15A1E178F22D96C4EC22E90EB07EC066CE4A19BDCD66D03CAC9DD906D9D85C630A7E10F118D83DC7618AFECF90F3CD32D265253A05FEACD7DA610FC868BCF54F0053BB7625CE2E2C35C8A24BC8F3DC294F60DF8F345ACF03B2D8BE69B36E51B49492E8891FC09787527B3BEB02E6B2B69158448AE4507FBED5C3FEB923854656B642CBE0176DEE52B92EAF411B5E1480738476037D52D7AC9C04D909EB7AF11D98BFC66DFFE81F19CE1AAF2E3C646679B834CE0030A6E3AC7BE93027D2D7347B9165F9DEB26CD54F33A90A3AD5FFC88044202208C3D1C97B9668542D6F1DC4E1FD2DB6489392E9ED43FA989E5CCD6CC63E357D516167691AF5558541513B38D8DA32D19133EDF12E1D161C5873BB423B4E52D6B34E97875186D0DF7BB4EF4D05023B19274FB1DF47631F6282A45FDA95A07F8D5B0B0F814AE31CF30947FFA65D940C88CC191B3DD031897F8647D0F8D68C2FB79050F90EDA905673B206E6BDC844875101AED46513041695E9EF151B06AF764BBCCA82B0C93B9D26AB96877B49C9368C972E5D42E2CD41B3F7AB17F8F0B3EB1D0C284C699D9F5523D6C5E2F1E33747E49EB675CCF1B68D2CCDF4C7CAFBD6B1254C141001BDA1E8A9FF6F05C8B914182BC4348655D69D7DE203ABB70242AD8851369AF610CAC22E62A9B300F53ED948BF17D811B6C6B65F2E858E645F95A7F2DD7A9A6D6C2D627BDDA4C852C2AF523F9D03109335639009697FF25A1C67E3100083BD6A741A5B4C8D5567A85820E3D9CC6A7F03A1B7C902C75EF1DC49566A0E3A12671097F086CA024E61DE92F15303B0D6613EDF5FF80A5AF17FE2613437263899D8F66DD19B34A7887B72F416B8DFF7498EE37590DE4B1AA099E9AFE8B78D139238AB3473B60BCC70616F6ADEA0CE912C640D4672C4D68F2DB405ADB6643D7C82EF4F4C95DCE932DC8C96C870B1B7C0B91CF5150EEEBE6973068A3E60C5DE142C96A2DF5495E1CC3B3823608116D0838A5DA3A8AEB40887C08E58A62EA753FA3DDD0BB615646CC2A5B185C7B55A7DDFA9704C4FA0A74A2B1BD579C24AD9110B103A6042DC329CBFC728152533A41C3DD19C7F07F5DE5C863C97DA162E01FAB8E70DC91996897C68A173610B61558F298EF0A540BD762754DABD89B89334A2F95A9861879E0D23DFCA4DB8F04DB6A7E6A3D67";
    verif_kats[2].expected_RES = "9C5EFBD8FC4BC59259C5528538F9546FC47C6ADA017628AD039E841F3EEB41078CFEAFE6BCA288F8A1DBC40A0A8DD61D7CA0C5DCD435267B4352CA2E2F3BD346";

    // Iterate through KATs and validate
    foreach (verif_kats[i]) begin
      parse_hex_to_array(verif_kats[i].MSG, kat_MSG);
      parse_hex_to_array(verif_kats[i].SIG, kat_SIG);
      parse_hex_to_array(verif_kats[i].PK, kat_PK);
      parse_hex_to_array(verif_kats[i].expected_RES, VERIFY_RES);

      `uvm_info("KAT", $sformatf("Running verification KAT %0d", i), UVM_LOW);

      // Writing the PK into the MLDSA_PUBKEY register array
      for (int j = 0; j < reg_model.MLDSA_PUBKEY.m_mem.get_size(); j++) begin
        reg_model.MLDSA_PUBKEY.m_mem.write(status, j, kat_PK[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
            `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_PUBKEY[%0d]", j));
        end else begin
            `uvm_info("REG_WRITE", $sformatf("MLDSA_PUBKEY[%0d] written with %0h", j, kat_PK[j]), UVM_LOW);
        end
      end

      // Write MSG to MLDSA_MSG registers
      foreach (reg_model.MLDSA_MSG[j]) begin
        reg_model.MLDSA_MSG[j].write(status, kat_MSG[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLDSA_MSG[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLDSA_MSG[%0d]: %h", j, kat_MSG[j]), UVM_LOW);
        end
      end

      // Writing the SIGNATURE into the MLDSA_SIGNATURE register array
      for (int j = 0; j < reg_model.MLDSA_SIGNATURE.m_mem.get_size(); j++) begin
        reg_model.MLDSA_SIGNATURE.m_mem.write(status, j, kat_SIG[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
            `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_SIGNATURE[%0d]", j));
        end else begin
            `uvm_info("REG_WRITE", $sformatf("MLDSA_SIGNATURE[%0d] written with %0h", j, kat_SIG[j]), UVM_LOW);
        end
      end
      
      data = 'h0000_0003; // Perform verification operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h", data), UVM_LOW);
      end

      valid = 0;
      while(!valid) begin
        reg_model.MLDSA_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLDSA_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLDSA_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end

      // Reading MLDSA_VERIFY_RES register
      foreach (reg_model.MLDSA_VERIFY_RES[j]) begin
        reg_model.MLDSA_VERIFY_RES[j].read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLDSA_VERIFY_RES[%0d]", j));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLDSA_VERIFY_RES[%0d]: %0h", j, data), UVM_LOW);
        end

        if (data !== VERIFY_RES[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("SIG mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, SIG[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("SIG match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end

      
      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end


    `uvm_info("KAT", $sformatf("signing KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



