//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the environment package.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
  localparam bit     AHB_REQ = 1'b1;
  localparam bit NOT_AHB_REQ = 1'b0;

  // pragma uvmf custom additional begin
  // pragma uvmf custom additional end

