typedef uvm_sequencer#(mem_txn) mem_sequencer;