//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef struct {
  string SEED;         // Input SEED
  string expected_PK;  // Expected Public Key
  string expected_SK;  // Expected Secret Key
} keygen_kat_t;

class ML_DSA_keygen_KATs_sequence extends mldsa_bench_sequence_base;

  `uvm_object_utils(ML_DSA_keygen_KATs_sequence);

    
    // KAT arrays
  keygen_kat_t keygen_kats[];
  bit [31:0] kat_SEED [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    keygen_kats = new[3];
    kat_SEED = new[8];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // KeyGen KATs
    keygen_kats[0].SEED = "38359FBCD79582CFFE609E137EE2EFE8A8DBCBAD18BA92BB433AB4F09B49299D";
    keygen_kats[0].expected_PK = "6924BB4257A7B9AFF095C30BB35C6AE4198263120F8039AA4E78E174A786CE008301E666F59D3EC5044DE456788FDE19EB39677B5F9FE14150DA463A706F3BAF715B95336B2D685A7CD7880713E4587BF7D857BF7E315696B8D0D9D49E142918BF0974E7F43237D4BE3AD394599E3D39BB7649932553447E5D5ACC3499930176ECD3A844A425F50D0511C9226C4B9A24F2A011CD88D32308E0312A0C87CC34A995823C65F4F0F98E50C37788CE38DC28FB8B9BFAAFA904B541EE712F6A041E0611374F6BF17EAC0BD56F3B6BF336DA9242070C2469A20C4D1616149A6159252011D299F93F986D875DD30B38A22549174570138C2BB3AA9CBEA91974F3D89BF5AE32BE9E58B854A2F8E86FF76780C03490F467DB0651C20B1DF60EB97A3C99D9BD664BE6A5E4C8A8AD4CC36390D7004E4BB421DAED654C357DA4D68498933EC71777AD64C2AE013C73EB457C68EF9A745ADEEB4FDFC879E774D03FAF6B14AAB10752E24B52D0F2D94D540A1EBE10F597E514442D6C13C2E2498E8AF3017C52DB233A90717DF25B4D072B7D88EE8731D16824C95D1FB983C449DEB466276060FEE4C7EE381451F232C29C7C3220850C61D1C3C00DB1CD9726A02A56609F3A65D3D164604588CD9B431412F1ADD914C5C2DABBC90467C0C4EA5F76E24AA618765F8B0636D7B065E1F4E6F622EAE17152458C766586772D363FA99214F472B0DB8A1E49D82D0278F2958B0AAA1586DB134BDFD2438742495007E2FE5B60E246399226947A12EA17631CAA534687CB75C060B4797EAB8277CC4F8A7A20387606EFE2DBD3E736249277D90FCAB992A8C99E85AB03EB4CAC5D88553958528AF92974718135F1D0C793EB000EA0AEC3EC1858FDD18688D1DA27278DEBF2CA8110BA4A204F7930E1C8CEECAFB73F75DDB34C5C55968A7933058426B55D039F7292AC43F64584F6DF187A1D6B003F514CC13B26C2F348195AA321DE6A27EC11348DE50D825A2964C631992E4B0B425B1BEB4F9600E3ADC4431CF2E88B4223D2DB663C3CE70EF85DDD56A9BAF138A9D7EDD894131C3A8F41A04EF9F86752B72181FABB37C86B877E61D60EED95EEFFABE6376E14ACA817C5F41961AF8A7849BAC094917B2D132276B6B3486AFF950D23D4AADC24CE98A5269E1C69917960A31EE09A527C358175CAA0CB1B018E9526D93534EADBACB52B273D735E22DD0D5C28FA3E47CFE90B5215AE24F146C3464BFEAF01D28DAA553C1E94428A104A9D78AEC762591E8879F76851CFB4648566721B0CAC1F14FE16149A9D8210CC8F2F50DEF7B46C843BE93BD8D55602493350AB560EA5BA17716423BE0EB8360AB109D8FB18BFEA040847B7335145D4F200D19CF6FE7BAC917F426C9B3D39A9CA4329818F240E7DA382761072F4A6505EA8E76C1E446FEB6625E38DDBCD3CDA81E83BF768F3E01D9D263B367303AE156C0B7183364A1E7941A09298A3ADF7BD231E6114B9DCE7952B113F78163138B9266F843F1ED97D9C2B163A6E8BD4C1AB4E179367C5AC96CECF5050FE821FDFA44E9E680B61C6018932DF717811459AF2542E2CDE77178C2E9880F011E405EAFA59C8CBBED76E5A1941104B1B9D3A60491C954755E02E894103F1F4977475E9EA36609FD67C9DE318EDA2370DCCDBB9CEF7AE6360905EC220838C9769823441CDD0DA8EF0ABE5F2D1D76E2FE08FEF53DE1D6166AB1A92B1AC093E5ABF7658C4B57287F2D1FD7B82DEDAF8D5A4FBAC4B35D58231694E162497578ABD7AA7C8FE7B3541A7F18E54E8B7F08764C5E68449DF655901549832D628FA63D2B2C5A150933994A9863317AD40D778D9D2C05C7898850B90173223C7A0AF890FD7E66221B6F06318B2ED5E199CB424885AB841E7A4726FABA2F9BB53BC3236434C35FBBE4B1A0F93F50C37896C29F8E302AD31ED3331D620E3B629455101A1F1CC7BA5E46E68ED4A8CCC87B4DC75BC0162B6330F833FBA2575DFAF5B5F28BC54FF2BA81E7A47313C15482B605E66BB38C6198F1392104080FBE78B86B1BC9A6FB881F5C7820147E6BA14B81ACCF20CAE96641094C216902EA5C125F6C935A150D7C9ACC5D9E2E5D90E38C0503AA9426017C76AAFCD5261B506274EC13A9679FB09796027A4BB759D928279B94D841A097393BF7E5BD69A496CC3DECD2B0F07F83392AADE33DC51B2A84F6A07635DC0EF57A9AD5959B6A50B7BA509AD5B11FAD26B419F9F1E3F9C7329B5A953D7CC87B2DE210611CF52A639EF2B3908012CB88E1D6F57625079CB103D6C98101A11BD2233B65602CA3049BD320520419F76B061E3598DE38152C88767D1A24FBD02BB10C38EACAE317DE6BB287B4D2CAE5DA0214965D8773778626E9B972859D8482B8D0547E4F56DFF87681D5BC5120F613FBBD91E1F14E6DEFE672E2A7EABCBBB9B11082C5E700AA0B1F7C1785FCED19A93AFE7C59FA2519BCDEB494C3D13B2125F385323B816C68F8F5628C7C2ABFD0278A337073DA74D16099698C4B114E8A8CE344E0A15D0FC7ED497B001D53D4C96DC3954D3B4B956CB9D2A272C51F1559B22904B40CC8531E40CC412C68CB6EEA4A4090B38E2797329985467E818A524D3228EACAE7825D3DAD2EAA422FDC77AED71A205DA7838D945E7FEC37E4DCA67E504CE35E5B045F56F1E8D7529EBD6F1AF7B6E939E2B7AB4027D37A5135D172DA1AF9CA2F728A6F37DE60DD23D97D11E75AB1FD51F8E9A1397E5822159DB583802B32EEBB4567ECE3746D1AE33314785643DD2A0741E7F1BF2D261F22124E8DDD08C640A48B54717517C21CD325328BC239CA028B2630D063C8CC20BE9BDB48502DADDE73FFED5963816533E020AED1208536255B1CCE985433127FF4F04D5B1E2F2108704B8B966588C0156AFC2AE192986FBEC443BAEF6CB85A6F29C7792405A24114710AE1C746444FDF5FB659E5E346826207B8C54463A0617CE17FF33E40F931FE576715C932EF29FD76B04A69B58E0303D8EF25678C8B70AF12E9045591C04E8B77106940415177E868593A09C7E14619A4B332F9ADC3A658B86017F32656C5429C115E110037A8CC7E544677D2DD239A59D54D0F3C7460EC15208346BA56DF5086C5DBCC41E0C95FCB6861C2C0C32AAF3454EFEE2FFBA214B430EF248A59B32444D8D0D3DB87C9D4B1536D157728EE7585EF532776A003A023C0AB0E9FF557108C390684D565A665063266AE6670ED53B0FAF8FF67829BB737825B153A9338CBE3DF1A462849B93A81F84ED07BE6D6240003274737F618DCB26E48252CE4204DD3139FF6876F43B305D835620FEDF79AA67433DC25287320E9917967B70B2D866D17B698BFFF2B3AB9514949E58B57C68A45412C1FC421C768BF5EE8A10C8AEF56926F51EC62C11569F31AA517868E5CAD89E958066EB9EDD7271B31CB4B1D6CE211225AEB5B57F749719DA07ECBEFE03881DDE3D81E4135F2DC81AF779776C1B8057162A6C982FBB4DA6A9AD284AB10C70022044F46D400BF6AD7182D197789983BE99227979A1334BA149D869BA1C4088123435BF978541356DAF171F33ADB1C97907A0FB5845074A85D26F546135AED0F91BE4539C12BF9411E4B556F687D069DB6B21FE2B7F321887448CEA55DB19FBB8B0482A55AEC16738D74CD265093836BE99D4FB53E9B014B037CDBFE9";
    keygen_kats[0].expected_SK = "6924BB4257A7B9AFF095C30BB35C6AE4198263120F8039AA4E78E174A786CE003B9AC2C1422A1AE802DDD7464D3F32729A3C7DE894D506ACAD25CEB372EA3149C98780DCD1314BAA29B9B807754C47DE5DCA954064F28528B815FE27B79AC506B3AD7629D2C971AB8F282E0C6E7E5548EE0E113242B7A0E064A6DBCE30C5619B19800889A04404B50013C088C1302962124CD3B4910A352C43123119996522185202C38523440D90244A1A30224428618106291897680A200908326A44A44C4490218A16689AA8511AA52C62468D04C340D3862860A46013187084948C63C04404A92820082043162A23292D1AB12948B60921883100C53000C48CD98268E1304C6332450C328618083191980D10B8709B302264040893A48C21C9700C35715B000D143122CC98102104809B28641C308021307118335024254408178CC00848844490489830CA440009195119230C52200E4906321C154E194885132549A3000408156D20410CDA4252C1348C00316943822464946D1C81110196214B0200CA2884CC466451186A181000A4982160B06803946C94485180404692222C23446998264D1C01085202208AA6080A316193400E9CC81181322E21158484C24100227254226258069248484411270404C011928245A1C68CE33266C138725A86010CC99084340858A86080C070D026629B302A04296904108D0BB904504628504824D04805A24802C3208CA014004138214B240104B5494200000C2428124084A220449B069063C0888C14214912105416242087445010850CB564DB2441D042299A168A21B44C13B77010C085190269CC40611C4846980625601446E4226224272262242944C62D08318420322104B4610A3812D92844A40820CCA8290B21310A3429032140C1A26C8A161252A664A3B251042951C4049163B02D1444308C40660C400C01A52C09942D62C61103985019104D19A828D38640C0306554A671E0B4859B8610043669D0462918A371402249004385CB4028893666412269A42851D98029140721DA80911B26505BA0609942715088491023095A902122278E43B2700CC94CA402709240100A397002360E113041D8402D1B246DC392614C868D21B800D3242212C82112998509160C5AA22409344210A22403428CC0B28D12B66963340DCCB065A112114A3869CC148158440954A6800CA805C4388A8406019B322D831290090260A1288858104124400219344818A04D001062132250E338219A962153088051260199C4281BB97104978404052CA0C210D3428181424D61846C5A30491BC224C02028CA922D4A90100427864C962109194514822C11A69113B80403187001A2515214495A0230CB302C94102C00498609A025C2124C1B026940A444411662022528DCA22D0016425830665B8624D42448DB260C4C088501904921244154068402434A244205401448CA4484C0420C9826049CA205D1C2511301861CA150D902500C39868C0031220548D31081124805D1086962382C0A23709B4472E3486E22967014336CD8902903004963208A039125088921C0820C994032C2344E4B9869098044E4046994200999246D09A96001292DC842288A3402E408700C236E0A054964442A82C800024831CB90501C056812122CD0800C594861CBA6099CC08142B80024418A94204042144D19466218050924336AD400611248328A047293B46962C27141A68944963162304683426C00192209464D8B0649E1B070424431C180659C002411A83113212C4B46281B180D884270D1B00D90C845DAC248591426224400C2944150C804180000CBA62419021010890C18222162A881C89248D3942082067209A8900C498A41862819C5809A184D14102E2212520008120C334563C63010934C60C631DC400E98825060022AD22240E4062DDB320ECA324ED4182408C3284AC268E28040A1C86451C265CB166023094C820468D9222E1C499242242100370EC812726408250A202A58240459164C08173000460512904003072152C0641C836D9C322E11158A1035885AA08DD9804803B64C0110651086401101420AC164DB224D64B25102360D93463114B668638429C8102494300819370214824588284054A8299014126136120B098CA49828C292454C006063C481C03625CA882D244030D3A82DC9C825D2844800329250A271D3440D223460121312868C5F8620794A050E20D0E1011786240EA664F2F69BB1B7E30EC66B1A4A0BE59B79F2198AD9804483E475E53B3C49CB0CE5EF92912AF440F23B995813D11B59F798E93C9D13539817C7AC68CAD1AA1AC27656BD0C4797E9C8EC17784C1A327A9DFEAF4D6191EECDAFE049B733FE39D5EB4000936FEEFCF82928E9F94CFD5CF4C1E3DEB1433A47F6D328B5E83DD156D0182DC692347591AA6F732CFBE982935FD1846CACF4CB8515C55AB85EE5AD44CB09D3269E2E6D11780961FD131D5E6FBF89849F47F2B71D8283FF25385E52B07DBB266C674CEE3D0B5DF5A56D8BDCDCFAAEE6A248E71DB1345AFC597CA830A1A35B4396EF4C1ADF9ED01BCE9B6EB637FA24AA160B9076BAE30559F8B29DEDB3D25B79064AB0CF8B8D70ADDDEB8B174248D5AEA4D18DE43B8938CDD2ACBA5477BD4AACC3CE595E5D269FE675210D23152B04710F368428794A75F49B683ED20DD647515777955A8CB38A36AFCD2CE0ACEC4F0DFE807702D1EB3BDE72E9E085AA4E09EB1B0947413852EC3C0AC52F06CB959C85394EB3748119EDBE6C80D2D8F792CE0D915E4F4B151EFB135E7F4DC97D858141C57F70417B43A6A126956978D78EFB9F037243B4CB41DF968B7EE5B52087F05AA9FE487BD16C0347CF1335760BD2398AD54DDA00A5AAC446D80B1C7998C602192ADAFCB809D14EE328641BA3AA00F8D29C3A848ACBDC1946BC0D35E0BE0F8F7E3DA3F68D9FA9768F5CF275534A0ECA9E60FCEA38F1E042C316143A767B33ACCAD8C8D66C70C75FD1F0B2586B653AD4AF54E56EF06933EAD31DE365D110B9C4A2A98BCBA165CAFE386F887C72156EB14FF0DAD665616CE3CE65C1904F2C1747B2EC2B5C9D6776BCD79E5AC64B7933BDDEDEDDBBC725BFDBCCDE2FB375AE2BE3537BDF89BF4C25F83A49D6A6A8D0761CF39D620C53ED837D198255CF5B910A6DB57877DF92D8BB6E9C526B8C4EC93100DEE0500A210C984583E1538160EDAC2C6F866E7F5D99D7B1B81582F5D0EBBF2786E3F556013BA9B6F656EB798838EA0579201A95D56BBC3BCDB9511AFBD4D81288896F87108C077F1A81A3BD297BB124A80086890242995E03CF42A0C21E272A9AFA1DC103463D2AB494F7D017686D31894DD2F6EBB0C3CB6223EC79C65D45C1B0D4EF1961F16D653FCF25977B651EC51A13AE8D4A3472EE71969A7A936F5DBBB9396A46D97642358CAF4894C9A6DF84A59C5962A6990A76F0614890169F001870D49CF2E75008CC4A5D85E72DE2D6CF3FA71852253522FE8B0E423CB417A38EB78C8763C3720C04E67FF88979EBA09E34538BB523B99B8E34167412F77AEA894D83ACF946FC054D0AF47295E51ED83F7486940A4D41C04AD7EBEE610BF1D03FA54071D51A1509E4F49163A25081BE8790D087F5F4F05C88550FCA9BF99C9BE5953D51DD0845C93E41EEEF62E0794B2927C4F5ED9BD3E34EA9200A79DDEB4B2D8F305FE05F827C7E2ED186341CB5D1152FC80104E0E13683D941294C778417164B684A976E56E78DA4D17C3C73229314870B85C455C23B830B9A28A3D8C0B566426DC169F326ABCE2EFFF39E9B199AE5C1292B6F2EF37AF1DEA9272C8D5423DF8A5632F991E14DCA2514788B62BE164828E9ACB893DDA602A5E2FB9EFCBEFD95ABFB82D2B02D49CC53084A49AB1BEC23E5B4C8E714CB03405F1BCF7E11BB59729DDC0B7BEFB291276DCEDACAAD39A2F01C7DC98B9E065EAFED1CC8CE3E848080A2FC5B98C9F6BF5040273342F0312F8B9844594A503DD3E6AF1C9E35C1032A4A8A5E7BF33A82F35E16EDF8C60C90021D8C0BA4C386245DFEF09448431D8C00D1E26EE4D8C77DAA1A705ED4792ACB4EA27C1566FB56683C43BF67842E67534CB3F9677C8AB9D0EEE7827CDEFC223AC948B880B5F1CE9537272932002C1A4DD218F527166EBFB2B2FA2BF37246ECDFDFA72B6DA11C30D1C7D248AD64818F691D59B755DAF71BED9AB5FB52E03622A900D66B4C6384169BDF9EB61C02DF45FB76B1A26F34E938B190861745C021FA876200C7FC8E222DDBFAD8BE781B185424AAAFC65862DB132BEC6D18837A1F58A876C99E63F51420B83F459675612F7ACF80B4EB1DD0721CAA1B4970DA608679C6383E817FE16B66B19181EDFC39270C7E917B1F10EB7A011997E967853B78E00CFD58D224D933CC5A995532DCD4E532E4030515F4A05B331D575DDAC29BAB069F09AF0D173373DB1EC2B6366BB371008A2386FD88BE77F5ED5E198CBE88DF24BC6E393FEBC10C470A72D47C0F834653C9AE800E893C6BA68EA28A838FCBB69C3E964A5FAFC2067DD406B257C98DD3979EC7C7ECBE96A33D85515DA2CB6AA5E1FFF204AF62DD4119A0E48C04A3F2B38660F52964D8D4AEE146A9C53C31906DAD0FD90B5D83B3E31B690A4C4935249981BE1F1A85EC6E0FEE4C88F2D89E2969AB8CBBEB501916558D29EA7C3ECF1C9EF1A04350633B4CDA737DFB151CB5E7361173F3AEDDDF527D73F2F9D5B6213AA68F883E9A2633785EC6BE642A9FD0F21A42F6B9DAABDCD1E6ADBEF64841B59686EAE3EC88EEF0A9CBC12BC012622DF2DD93A86229044AF2F260D2183F51E833EE92D98F0251E3F85FAB74CE367B8B7AA63D3CF8C8BF4D78358BAE0A0241E210AC69353087CC7331357EB4450F9509CFE595F54032EE057754A8EDD746CB9282E768DC6B830C5B4A219343AD124EDB3BBC42505566A7038C959BC35585B6055F1968DA243F778F4E46DB462ABEB93B81243C31EB59622EDF81F06CCC61D2A6EA73E109C387915F277BCF1FC11105BBA70293C0FAB5C065F23BAA19290A302F08091107A4B1D568852622098383427760EF8F2928625BDDA5F514C5ADE959891EF2959F248A3532BF9D30E714059EBDEC958708F8A83C268BEF2682D603CA886347E198FD68233999C77D30D7455DE6BCFD0144277062B304BEF0E34C5A9D8D780D29EC2321E07340771C46360483ADCAF12D5B79FDBFE2856ACE8859F6B12414B3F7E8BB5813498960F34FDC64FC848579CAF9DCCF19B4FB825ED5716DCCCD6872CBDE3831D67384942CD8A9EC4BBFEF5706B8F9F05FE1E8FE69D3EA6A8621C22144177B1C1259E1A79DFDF89728887BEF1A70482556831B672440E13FE3E3FC8204A02EA1EFF19D95253887285BFBEA16A0F219EFBCEC30A8AE86589A5703103A8A393FA6F6B657704AC677C14CD10D3D62D13FBD378C2DDA325B61B85952D51293871E1FCDC948C77BEAE9A6F0E87CE1A8051C8F8087685C12624BDF58380ED66F55B43DDD6D362173A5BD389859C17D95ECE3AB732639FFE451CD103EE4854DB2F39614F658BAA384BC9948D0714EB48A887143E7A1FA4B690C22B492A70C612B59FFD2D6B3B5E99C2003E2C359B1E62DCB620C7A246A7B9B3246131556F2F3D513A23C6A9FD2280ED686D767CCD01754EB4C99692F2B380C36081344C1D35EE1949736B6976F4852CFBE64FABCF11B9AFB828576B4F9787AA7D03E84598A7143EF7311FAF2970E23ED4C173F985D6450165AE3E241A18234E74FF3DDB921A5300B1C4FB6E432E698F53F66E38C07BCD6E77605DF4624D579076292DE1CE6FC6F0081A38BD92D39B24B73BAC1C52BD68E9181D3DCD0AC7534DB48901E5984F9902557BFA231B2EA28C3183262A1B2221F7426EA88A5816093A5CAE2CD5D59A9390FC93A2956944B064CF013BCDB67FB423D1328D2C6D7BA329013FA2D30EFD69FDCA1A95EA6D06C7363534B2F3F7DAAFA296EAA09B3668E9CF82D9BA959B32F3CAD3C10C6EA48611554539C37DF6BCA3385EAD3FCFF96D372B42393B73C8DAAAA31506EE0527B7FB3E593DCCCA57C8FBBD4A3C7F8A53899869132FBC3E4050607BBFE29C675E3945E74A31CD531BA7AEB2E2F0CD990B8F983A90DFEA0568F0677EA9563F7C479DE968940CF242992692865CFDA89FA078BBEF49CE4575BDFB380366011C8435F12B42D9AB99AB6A31912C4354149D723101D1365A65E7CC68D82E30517773902FB38DDA2B324E7208E987ED287D092E7662A430241BFCA552D314127E38C8597A89519D4F1E62A79465AD5F4EAA3FA77CD98326D2F92CE9852055CECCF62D63CB9D7F198AE085E4D45C8E48FCFFE593AD652D9154167BF3E6195810A445AE158F1F9A6793363AFC1F22CA882FEED3A5F5727CA76477C5F23F0FC8700CDC6A5BCB2B20B4F9266351D304A96A82BF5F314AF685C1C707C92E3E847B7047D689C70B25E5501CAEC9919626F4A0FC81586AF1EC88889B423387D5D95482618A650E80B53B07CACE3228940602E3DB47466CE9BCCB6E4D8AA61C8912583E810B3B2E7E9CB48BD403ECF08D28C70AE0B620859C1F09B61131404C3D5BFFCD860E0F42AB299006230B2876D77DDA91C8C62BD93A844E4B344E3255EEA531C6C458D04ABDB0FAEF2D1C0B4C55F570A5A51023F4D4EFFF59F9ABE17922FE732CA71BCD434AD7710B84CD4AC9F2507A06826562AD7F647826F9DBBE4EDD23F124369DB8526FC2B4D52F0741415F972BEF6A935BD812A56C8221B7DEF0F5106BC01E913E3D43DB86C2BB4C7E0762663C6DE788721C2AA07F8954887E2142F2E914A099EFC0AEE1339210D3E53DA3ECF88624B1119BE34010B886C80F51D1850838F2150E72B042AF32899C0D3D7B02A57F8CF263A369562E4E945A31282A502A95EE9BB0316C6861006DAC17F936F54C4C7";

    keygen_kats[1].SEED = "29B4987C62218C19C77D695EB904AFFAA1BFEF6A52F138604CDAB1534E66DC10";
    keygen_kats[1].expected_PK = "4E130489218BC6CD1A9DF06B2586365F4362D8A007563DD1BF7D77F29663CB459F1B080DCCA1E39FA04CC66B9DCD4A6CDD2FDC25B96E87D778C068A41D7D4AB8FFA0E156AEF370568021A0F56EC60853AA4579F7C7151A31A7A8E5257D791D06ED11CB264B658467E82EC5EFEEB6FA224577EEB84D4453C82D821B87771FE57B10526B6B003E94F9CC812731C08A4B9FFCE90A06AD3134BDA3CF4E7E46DA7BC775B95116E96B53817CDA3FD3BC4D6F612C52BC2EEEE4153159B6D223E7A7B20EAF926C822DD064375FD26CEE2DA8DBA4665409D5A4F38BA2464D393FA00258379038331E4FCE0115988C634A95656888EB26E95049435440F42006C3515C7BCF4EBD138792B163ED11ECB45719D9B7821D6F7768B631D67DC614CF595C42FD2255252152C38190A5E41BC5868839EFD2E12DD73AFB61E8719C0ABC10679249DA931B4BBA405A46C3C112A4004A8E3A273965DB3AEBD8CA5D2BD12584160CB21369B1C5163D111DDBFC040CECDAE8B580B038B0D476211B05414A04B72AEA2FF2BE302422CA22F77CC5E4B576BDB838FBCDE65606F841030C2EBEB821619EE7C3C60C82BCBC3D55B0150A72A95EB2363121B925414138674A0619E128EC73EE4A9868D257F79F27658657CB72D9987FD03826C38DE6509F97B25144E4D0FAB4F40A3C152CCEDD908C50F8EB12E775CF512337BE1DB1AE9B320541EFC0DBC70ADC7C50494295C11D5770D6AECEAE9EEDDA468AE90800474D80B5BAA4CFDFA0A56F3C120C8A2397F31C429F915D1E748539C2A60BF05FA043E93D503FFFFD538D5B22BC0FE8498DCF20EDEBFB9FB973CB00EFFB3B65DE718292D783A16BF01301AD2EE546D48C0F44A05323EB15137C0527CB1A55775A6BE5B0F3862BD8EDDB3CD54F9AFABC42916DB1473DCDF9FB115A64F8EE011F2CA6D11528384B3757711ACA40979C23E65DF41F8D4B2D593C1351B713AF8421970D9ACD3F7E7ABFC764B8CD985159A78205F20C7A478CD987A18325F20D30C33B172E94A7C8F3B097A0627EFB6DDF787973F4B410EBF38E3215B59A4C218FCB5973A378D9A2CEE29986A61B841069BAC816147D0D8DB1BFC8E7E0FE811B589484F19FFD03890861703A27A0C9D451048C925C40C888410044F7420FC25B6B79F99E1055BE964968C354C917F3F981F7B67D1AB451E127CB50E5A1B8C3F179C3FF2175DE548D1137297555BE12489E6F3CF2831DD0E45F2E4151011DBCFB8D55AB280C0F0B5A81B492A33C674BE15221A990B800D9CD5DA9048FDB938633A3BA965398D8FF1AB77F301ADF74FB7AF818E4ECF587416D1CF1BD0F50A65D5EE7EE34E1B6388A3FFF8063B12551BE96AD882EA8D4DEBD9E7DEB05990221114784E7D1092FC01F7BEE9EABD72D3F49E572BF79C771F3E912935C2C71F61BF53EEED86D4FE1D85D702E0CD0D322A92C39935C9ECDC838242C3C97B708A40CC8311F72127FA66F6B63F640C1499F1C70AF48179629E404ABDD56518268BDF1B55F3A6A61E4836B881CFE7B64A9663402FF2DDA2997BE6A557580477ADDC419D5932324306F4BBD3E014CDD8D8FC9102D1431BD895B0809F8BF9214932E915FA0CD1A67A00DFBAC207189D9DCC0A5E1842B92233B8336F19868F29EBD31064EA8227E157942ECBB4C05D40926B4497F277394A7625DE21518C1CF3880F6E23A0A18918BC441A8E7A2E63DE4A37EC35E559FC5FB0CC0E016CC7FE06752866DFB1117B07B635663F39974FD138700545F6B64B2AE401EF894DE97FBCCD34ACBD5CA3AB9A63864E2B0B5B12306065268BF0427478CA944BCF25B2AD50BA6D6481AD0D40EADF2977F12D028421AFF4556B7C450BD8BEEBC697005FC656051E8EBEB7F288361DA5F91AED8F578DF23BB964C68107E0FD6B4C022779F84D78B31F2D152B07D1DA564D425484A0A5F223C4EDE705CAA2652179FBC9A65BA065039E2D531B80645FF9F54FB131F697FA80277B743F33588636A771CD9DDBD0511FAB5F1642A02E043AAC57618887534FBE5EFD1441028BA58D68A390A3DF8EBCBAE896170BAF3E352DB8C2857DD5EFA25E2695C157234115D136631CA96CACF71D6DAD9138B86366FF62C30064EF467ED753D8560E47EBAB157E5EFE8115907092BFC06DA6F33FF14AD29573D61EFB73651AB2B515E67E9215DDF86BC52D2DBF2A4206AEFC55411784D8A44291AC7EE56E9D124E1E69B0C5DC4E418D88D3AEEC568DC2CAB4D812B124C7CD91FA8613AB0A5CFCD6F668075DC4069AAA37DC3C7EA67C184E02B5BB33D604C983CCB9ECEE5D4B6AF74E6F44932937425B18438F3D5F358BDCA002F8E0596EF63BB934A91B0DBB69D9B3830A5CF6E1DFEC05629AEBF50F31D2EBBD9ED0894617878F1B9ED88F0F718D765CEF17A06DC288484062533681506E440A3C0E84C90119859C0978D612F0C062BE8FC5FEF3A4759C9E6193C66B56FCCFFBB6D44C713B748BD4C4A4FABB9DA38468CB4300437E5258C383EF438323F23CFC1D6C77304EAB8629A8910CDBB91C3B5C6EB81DABD2240B62E0D3C60C25554150F33387461C514A258DD2FBC1EE8E39DA5BAA6AB3E26AAD009EB78906B488E41ED03EFEDE7D7F8E67605D3C3131F4FE41C79F9C146B6BF51C56734BBE8961421DED7C16A44730093AE312563B6D98305DF2EA0527E797DCB46330690ADACA60C4A240CC42F770375EC7A49800FC573D94E168B053DE9B5B485A530BE485EE5291301D8A70F1FAAE35B49274BF0739E0E5DE495FFD791B6A3C5DB7D81BD7EBA6DD2D9E326DF27F2DC957943B5BCCCF7A616B41B2DCF2269B9AAC96CC06337FECCAD0A870F0DF3F1F1E99E45869ABD22282EE80603DACADC28288B4D3BCD5FDB39C176EE3E92592310B3A7D42B58AA477D832E113D696BDC4E2A5946410803F24203EE93C13BF380F4C84E2C62722F75851E54B0718FF23DFFC937BD3D1D2D787673E60BD218C102B572C874EE3F5971EF7F24EA5EF2A093B6813718E526806F270F7712117AD6BA1A91D1A3CA817F66B0F354BE66DA05A2EF3B9D05685C107C74E09EA8BBFDD182A1C7A6AB9191224E4BA13AF29076652B79419E11060A0BCC68EF8F97598888C12BA214AB25FFE68298A959B0CC755F00D6FF2688E20451728C51AC2FC96F53115591845AC9E330AED88A7387B5F73A136E598041F7E81BA18321A0E620F088A8A882C691E9D8F99E4C00AC849B3057069F9A5A0024E3015D613B773AEA1E1581AA57FFC246E5EAC3DA2A84A4E48B60BCFA9EC42686ED217469CDEC1912ECD07A5BAB69FE67BE98515D200022B408ACB03E2E927E3A77E4DFF29AAAE0D1DE55779FBE73FFD37FDCE0A3FEACB64DF225FA31324C3E276BCD4753A2594032FCD27256ED4F34DD2BA992C3AAEFCC89F89D9B46635321368F2DB71A3F9612BEFDB641A6B33DC3D8AA317476BC805959261426F7331DEAA84B8C6BD2142B3077BA40A9284B6DBE7D6C92DE0A99D0C1BA619946BFE2537BC7AA29BA4347AD4FF2F5EBB554E740E49744E3200B7562CAEBB9FF565990B6C79E917884F162973DA858811C0A8D2799F65AA7B3CC8AFEAB97204EAEB83EBFBC6A688E48E7FCCDFF21987AD436DF23C16E27F9715F7660884E553421292862B5CDB5A246B13E75F5677DB14EB5802441A3F01F";
    keygen_kats[1].expected_SK = "4E130489218BC6CD1A9DF06B2586365F4362D8A007563DD1BF7D77F29663CB45F5A174EAF47F9C8BB723ECAE888081EF19773FD058691588480FE23247C9886F403733B8A4D5923E737E3EC5A5BC019D015672BF421BDB6A830CE2F9D229B6D2275C41BB2F14A0B5632D21945070EE1653E97CC251C8CDFCF4068211CB6A24D68A1290123730C4B87141040164442E24B4251B05251A248C94166EE33450844251234085591286DC08915CB870C2326A2497109186095CB2101BB2485C445261344C591012D9286023950DC0266220C70100108413A869C2322942C62520202182948908153153166CCBA0000944501AA90412318851427254B66002222A209130182344931629C80689E1B82101426D52242C1C13855322229B22916290909244308A2861E0A4518B222813111218098100076A1921419302908824621832280C898CD434000A800C22238CC8981181046D13899048024E0386204342699C44650CC2895A882559A06812316C1127680A394648B651DC384882102DC2364A02A12C5BC02C24A50118912160A64D20219100164620400150321011A2808A360E94124C1A1525C2C88C43248CD0266109076498B401C1484E04A010620201DCB0818C066624170222151251327291800024272E2009450AB9101400668410260CA25000828198348854060E9B36321C87040093444A300DDB84899A484A1B474513805053B840A38431412429CBC248CB3646A1340E18A269C9926D48128E04183049C8448C92800A46450CA05102184D19150108B8315A060813446A5B48655494411001689A448800305012070152442CD83080C0A22581226A194500489250CB82851394484A1051C3046D89124D02922C2313400AB14CA3B4241B228AA012204C0401A144898C4271641226C8028A884600E10445C808699A00804A3001DB102618B40D0C3204DC8665D898499B140964844161862D10808510016C22000DE0A830C418044CC049923485C03671A3022103A16DE0207112A7640815208AA4044C164EA12066D98001233730C3182220460410346890B42454424444B89042C888DCC29090106D13464C98C66443048582362D620009D0962812C02C88B00C5BA805A2C8619A84694008321B87644228011BA74D081761D4228E82006A5A420E5CB86101B6055B32668800318010901BA631C0401101443010450111A728843426DC90648C306481300A1289681CB92122472E21482A242705E312401B994114808C4B40104C1681584488A24672D3021121444552425108172C4A902188120221A02841822D58224420C500E00030129844E04231D31226CA960D0B4909CC480181262613248D98182C18448CD39200A3C46888102223136423238081A22C582009DC90445A148EC93291E1463122C981A02462181384DBC285E100905A10655B262982B09180C600E0986059306D18190614276D0C24851110200429894B2288C01080A2160A48B08C62304EC0446D4114211C3392A102891C23260B1209D8340422C224D4368D041451539021E1C2608A841114132920B90D984292C4361203909093C84493009221156523257092106E14C3701AA470E146209096280B342D18078D1A373110831083102DA20470822010430860501610D1447288906DDA94245226281025000C334143A04993386624A75182082844C2300BC47121356D0A300EC24240D4024A80302591B860A3042291A08113940C883800D4B670801268620648D848064806602423509A346222433183A6210C04484130844994805838049324286300020CA485C9C05162B28499166D98108183B681C0340961B28541348044064AD8320941022D0A352C983664C288695208850AA01000A22D1C137001A50081928509838891347111222D43862CDB24728CC4645A288A1C826854B04191024003486824346D24336C5C266A8104280BA4501347911122280C4301192124503840CA20315A488A04B8509BC26421450DA1340C634072DA288224C28404006620B729E2A6258094250C4265521040C32882DA1286022586884690D9288C02403123A861C930711828688C0866C90206582088A4A445201560521832C092600A09519404042302219B0620D1C02801122D2089600AB604642051CCA42C51164C21110563C23188C20544444563144A6130888B3860A118904C3852EBFE4A5235C8D8FDACBF1F0546D7E244B119225B648A9D6F84949F1097FF2A302FFD636B8ADCA5B833657227F6432C2409C7BB078696CBF666B7BFA550E7DD1EDF40119D51EBEFA2862A773F05427480464D6279581BC7E8829DEF05EDAFEDBA3894960E2F9C2700C52EC53BA72C8467097E08805A4C23106F3559C1CCE2AA70C23DF45DEAAFA26500E17E93C2A9FA71062E3DD628EC4065F78E192CEE47AF2C01FDC3A495EF01FAAB25C9AEFE9431154CEDBCABA4D2E9793291F52F8AB834129044E3C69DA4F726CB6909DF7FFFD4B7B48C1DE143CCB63E84276CC00595C1DFDA1FF6B134DA457C2B66E893EB6561DE33F96F8426E0E2791A278286A6C5B5155AC2E3B90821828C3546E451945863C0E9E2853F7B44C296C454F991D091B65221C1324809A8F683DA113DE0FF641C9141D68B888E816602F165B46777F1157C4D6C4656A5E99BD0EE46F89047B0C4A509AB2C3BED7A175E45815C16F9065F49C7261959FA0F9CF4B6A5A5742AD6C4D768F7B7AF02E453DABE24AE382DD50458A1D20E4D9F30E98404061F927F26A5B6A677B2957FE4C973B42F2A1A9F61A7C4DBFC4FA590130EBE23E0921760EF05F25D6C7A61E2B0D636FB21537298EEB279D38FD4B85744CEE35D168590C53AC9AF082A1B0C7A46EBE5828C6B98BD89F562C1145DC5A54B4ED8F7997D0E48CF90D56B9569D3A4C4847769BA3D1ED526724ADFAB7229E5CECAB2D08E7FA9B096669D063CA3FD42D2153FEA0E703E23178233435AB81E7588C9BAE343FBFDBE77AEF158DBDCE8E1A4C3A69CDC67F3EA1D4C923118310930CD2B83BF534EBA764635D12E5FC86EBF2560D12DB4B24E4434C9135E4CB7631E0B8AD570C54584BA92B27B54A502FDF57896EEF6054D55E2B15769B53784C8D024EF9B10CF583D99CB4155BB4E3E9B2C28D382952C062F6319D26D7DCB0E946767D13B11CB870265BF829A93DE55E17AE7AC5D706CD0484E62DDE8DC2B16CFE5063EB8327460C516921C312F2C47BE9E71AF239EDC87FB8EB3F2D712609B615FA634CF9991DD10C1897654D5534A537A193741AEE36EA98D768349BE367F63E21EEC6D6A5086C7490E6F6AB0D7776CBA761A28FB5C3FB1DCBB4A5A90F6A8147C80D5254C8870725FEC69C93285A5A974917A7F3E6C7EA58416B814FDFED39AE3AB71A62B0CBB0427EA697DF596784EFD9D650990DFBFD2B5AED08AE76A243497ABAEC5591150616BBA7D7DDAE4D522067062D98FCDDEB0360C2099F13CFC66D001B18C4D1A8CAF7AB4C8F12D9E931F641AECD1F894BBBD3A62E7EC18CDC02C2580625B5334E32E565D4FD9CB7EDC25E9ED12D0DEFFE81E94F62AD696BD3F2BD17585E9E3D87AF16C9EECF24CF61F53669918666F8585A4E2BC34F6205F5DE856BFC767C4D0E2B67622416CCF8CB89A619B65D9B0D002D457C5388314DA854C4CA94EC466B97C8A55DC08C73F7FF0DA6D898B7A77062F9150E322FBE3339C62AA192DEAB57816A27EEA7C9BCA609E79AB10C88B0137811BCE51E17298487C287074A0D1FDB59813BB535AC57FA6DE8178C6CEBA4E6130063DCA5D7E256D173C11E31BC072BA6A70582B3146113DF433F93D74A2A72CF55482A1030DFA0C2C6A0AFDF5E9837D22F7CE89C9A4D81FAF4EEAC6262701B011CAABAD823B5CED6918627F66B1A07C3E5944D53E161AF56478F7598530BFAC4317BB363D4B2B04BC3D0CD938527437C2F88DAE1D447033A315EA49B2ECF62EC6BF95711A57B7B6C0AB04FD6706FC3553A7B726F30C06347F4CF35D989F57AD779DB038280BE50125B9A8AC1A2C84F9B8C7A650A3EA1533F575CA029709E943DD9E1F2ACE7757143A8CB9FBA11025D49CA9CECE240D1B63140C30CE7D0EB2311E5BD9CD7EAA3FE81E93607D14D5D329FD28FDB0E62FB87D448C3C1F85B42FAEE0DC60993EBCFA8D848903E55E2E987D34467400B8F50741EB573BB9FD41A0A5BA61EC07EBDB2675912DE28FECB52A40494245EA078A754C1B9641F4F2B6D7512944A83E8D1A70B7F3E62A13E9C456152F163BA359752A91A8F833373D6CA24EE0901657636FB2DA1E9E0C16A789ED447036002098B7D9D66EF633047792E9CB8C8CD45DA05EB5ED49377F060CB67CC33AD0D609741D0B3DF408F584D83910FDBCED95724714F4334E8C6AAFF680D5AD60C5A1402A97641DC8FA7B1531DEAFD369EFEA623F475694B04E8E5F52FAC99D8BA2D928E60C4D8AF2A68683FE7EE6D82021E35B895D57BF7F4BED6E2DE8B0D1DD0D0662068D4A9674AA65121489ABF8DEF5F2A9F1E2D36A8AAFF54C56E2E6217C7C9DB4B750207C5AA367A25401C7A3C7ADA45E1BF4E3D777D1306755FC0D69830F3BF262B83E727E5415992D6BDECD7EBC6DCE31FCB1EE0B54DDFAF20B522608870C9A0B1C9DA746DAA1E13A451FDD6192EE7E4514B8B99BAE4FA2107CEE404A7BA585FA7E1F1529E66DFC6435A1C26D3CF0CA13836F0B44E8947833F8DCD0DC2FA60C9E6303BB78E1C6E72A3615F9B3719E9F6A0D2F043DBC9AD7BFA803DA6FF03BA5B366B50EA314E42AEFAB8D2861462982115C2C7D6248EC74F7289A3151EEBD3DA0F43B89E9B5C50FBD0955DD803A3109EE451F96F5DBF1F9B42CA04724779F0FBE9D1C672F6BC478E919A07A486732817EC3741F231E9ED25715FB86EA804DC1B23BBF148E20DA21E6301EDAFF8813F5A97BD9F196E40BCCC824281F7C7F0F4A5D396BD2D3AC94A99B0BF24BD7888276A52543B0435091B4E94328164576AE7A572D2C4693DEED54F583D85C783BCD540A1240C40B68AD8DEEAA7255387029653228EC60AF145C2ECDD26A1D0B267695ACDDD490495CCC87BC1013C065357569790FC44001EFCAC9DD18BDF6EF505BF5C4FC555DCFB2A098108A1C06A3400C10248480C8B3836B26CE19BA22EE4C087C687559B6B6EFCBDA275926CF10F151DA7B2A0EC4DC214EAAAB6F93043437B32E0CE139EA665E2CBAFEBE56D6F1B98BC82FB299C381076BD1E1B0564F39FF03795794374269B3321C8E2E9BC6EE8D03084C3BF949E26B759E5A71CCBCE856FD0CE5FE7F0531178B2C80E2F913D777CDF265CA351FD1EEAF2650A2C8A52ADEFE7EFDA688556AC442D9D4EF43AFB177987831AD7ECA98C3042581F2389EBB972BB11C8D6845C8159FFFF7B2B7AD2E77F6FD4FE21E00A528F1C243D84B4793ECD4BE3F94E59B2B0435518B9BE6BD0633E310F254B822A66EAA384D7AC066C4F273254F3A2C00CFCC43C3A52FEFFB2B51CE1564A0CE3682727BBE58D9455533269FCE603C7F6872A6C07BB290C0B8AA95134D55B8D551AD77F071985EDE813578564EADA5632B9AE931EEB24D6966DC6863DD2DEAB2E3D0F4CB3AE862AFEF5B6D4C9288B1B3079C395924C67B03C415E7A8070A6839996C5BAC53E427A61A7EA100CC10F3ABF7D311845DCA174FFD06C3F05B88CD2FF32E9E44659D7E80F40EC56172C68BC5293820886BC47E8339CBBAD03383D099888E668AD95A905373D30CDDF91756C9C7C89F6DCD6E0BC9E9C4ED9A876F1568B49B6CCE9C520110BB205E307ABF68A8FEA783D1FF4BDE01F57A6B1224E9C83FBEA507BF14F77BC27BA0806D48F8A0FA1CC1DC0EEED7FEE5FCBEA5FB609D76413329F54685CEE7E4FDD309114F71F864A26F05A672315150823110947291991437C60902AE0767BBD42C57D6C97F5CCEC62207C8123E750945BA0BB444C894A98DB610ACC5703121CF8A93C7CA9CCDA90EA0938304651EB84D2534F2E67960064F81A41ACFE3560066DEDC1D7F954C01CEC3A8083975829149FFD8A54E3EAB95A076361EB7561EFAA8E678987F381F662B59A49579D9A2453AE756C133EB4460E72218696DF703DCE965AC32CD144C83819076D6D82D8B5451E0FBC384EA3A2C5675F2042F48D1D1A914B384DD0727CCFDF0A07218B3BA7BD10A55A550679C12244059D2DE9F76A4B1855733725EDB2981CF956D22223833FD43B9669BA21B38FE2C6BF49484BB4FE9E5CCD5F883E856DF05525D9E3BC452B73E6CB6DB583E3641D215019D0C48EAAC8C03D646CE537800AE96457CF187D3CD456D13AE4B657FACC6D9F78581F209E94CBD19B6768FBE0F558AB7E2D4938A0D2D92C6C8BCA7A01D7500286756E87C9A55F10BF60E23F7D6039E17CC6340445E297FBB213730455D0A7B33B852E4829D31BFE5DC6AF3CB5916176E4D125863A49592A306B9ED9CDBA4E2F40A4C8F3C85943C10BA10B688DDF847FA2212E374C64148BF6D1D856768696C6C8F04D213065A453530CA6964377687CCB2AF180ECA47260A493C8427CD418E91D38C50FA9ABF904E419A612881CD595821657C95729FDF8D1D965E80D8F8F82C6009A8BFEBA81ACF69503B873F92E557DCA50F87187BFDAE231D0164CA86E58025F51B0BCC8051D9A88313A619B87BAAF7B16EC52808CA8CF9856CB09A58B71FD67FDB4B3A0B88536DC3EE689101CC39F7F0418E3CEA104C62E83DA5631998DE88562499C4D18A98A1DEAB254C74334C325C11EDA989F98548674C19CA942AA95CEBBAC2A593BE1A1595B702B701DD42E89C8E65DFF6E104053815FE2D7D0908CC2698D2B6C26FE981025691A1680727A0D65C37B0D87EAE23CDA4E6EE98F7A981B9CF44B6B2752AD2337E02CEE156BF8968174FBF7EB0574BB62434D69EDE82D49BE6DADB3510026559B7";
    
    keygen_kats[2].SEED = "9B54B9C91E0201251489E07D1442A42D0BF32189D0C0CA8A2D4871DB25F531FF";
    keygen_kats[2].expected_PK = "9C17C88109B6927D423D887BC2FC24A5C4405C8E736C1C9D9A799C5CC09DAC3BE947BB391590EBCFB93BC00F569874F69780502C80C4EDC87DC9378294EC3D62F584E70AA18C0F1139DAE97590D0C89CF57803A26FD82F264F2CF2A184B2DA47F44E22306B95879CB3A036C918B6166E1408E59D35E2177F6CBD05EBE6F1230FED71A3CA9CA73F3333070A1DF3FFCBBFF32F82EE2ED47285D8F05809240ED1F91873D3D817AF74CAA85BF78EF02EE9B36FF3BEADFEFC436001A219770927C1756A8FCD265721CC8CCD367C7B19A40DBA1C9DEE9611863BED506F42203AEA72EF21026307AF0602437BD5A8E7B1B1F1DED44C4A009E785BD170BC98C839753F076BF7ACFCF3DB89FACDDBE5F5CDDFF76931C0966CD935102FA75A967C67222D5F8DDF2412F0CEDFA4C9FD94C6C58F26BA4954D872229BEA543107613C71994652F9268EBF81862CE4DA0D172233D358823229618803AE54608871866DCE80B988BC82F702A8C16C9A6E58B465C39197432152297524CCB00338067CC08DA6E2AAC288AA9B3AC40493A454ACC7786D6A2F261E86F4FC6A341896C2E1B7EB46AD1E4F35D970B5B4FF1AE8F514F6C78BF27A40EC941DEC16C95D9D91F869B578BF37E5164EE77DB6D38F7E65D9E703C6323750C24C6B41BCA787AD02208421D3DB8D7090FD3D154D9561B9638BC20BD55EABDFBD0F772D590EADA34FADD191F4FCD80C4B0A9EBE8A069270B89FDC2F0C54C5E9D835951E76E4255B9AD8DEA2092E806D7C62BCD7800E175C93420D7D8E3806F2B6F325171A80C34F0EC7AE7C48CF4664BF07675B8C617FB7944795070E7B47EA9BE7509BEC0514439E9DE57E4C6A2A64303176D1BC37632DE696CA7A3785943E299A1B152AC93D1FC8EBD3A451FE780098A13A72F4EFB4A41131549038C38815687150DA19FB3DD1CB611B9196135606169090D426B33C0B267CCB630172BBBAA67ED2817227DBE6FCDE76CFEA14A17A36B034977559C9E8AA525052CBCDCB66E3410DF8D321F3992B02C3CA8FEF477F2E22ACD2B31A89D194CCFCB4C41F8FAB34128EDFF327C80022CB9E15FD41ADEEE69F227CFFD706312AEE2C824FD281D62C31C98B2306D08A39DEE41BFD1CC702E55EA718A0C265E116BE6B87678927373592B6438B7FD490B2810132579BDDCA4FBBCC0764DD245F6D4DDB97943F52A0FCD190C71744C2E6352F4D0D2121ABAB3870994E21D617A96D77C195436B291ECD15E9CD29C6E05617526FCD8F853C8CEF29CEC0549073D4AFF72CB975D3B6F4EC0BB0CEBA04E35E69E702D5E1C671424EDD6A6835E0E9FC9FCD7FF16B90B039BC1B1295F88F724AFC6DF5F70C22A6E7CD16315F5B7DBABEE28B7651EB16293E2F4998A4F4640EA6EFB4C0E8F51B7DF809CD8F53A4C18F4F4EEBDB18F3CE2DD37F12E0931A46B296158A82D6F4980ED9FC9316BFD7C519688C0C4BD22DDE4EED750EA96898481D7790B95907F3D7E9323EC42B59342A52616E288717B8DE4D5550DE95560EF33FAEB2E2A4D9641FD0630F487DB670B9490D8F91F4E2E9DDB7B6B2ED9DABAE448622DC60A5F869C96E12F1B26A77B42FD6F513E9F8C0D53BCB5610EFBAE271B754C735787E9FFC5FE8778E967D713C2C3CFBBAF59B2262F1C4B8C0499EA77CD587A5296A819955781AC371C20E66471CAE28C6B098A6D25216F5CC3F52A258EFD3E22B010DFB5971B5EB004ADEB9D34375B157EBDFD3331B6A9D56D8DADA55AC152C3AE497A36269F44F3180C47EB8C315BC3F3A0C8AA1CC062C487BD917FC3988AA468C63856277620F576CD6B70BA66D3F9377CF20452DD3E7A8890FFCF309D7E5FDE1B2ADB2BB6E96ED3E8F2CD1F075D82599B92F74602A87FE5506E25E2307FA48D0C171E61BE15E10C3EE42398D078EB42049D44B0A343915F3A99547E2E27DA86B6D0B88F9529613412FF6D6AD459F30C1BBAD521E99869F1F01EE7540407D645A7B6ABF590DBF180A85076CF838D89F0BD53CA96759CCD3F11726257FF862A565217B82068BEA4BE94215F0DB4775558FC6D97B7D4F3254A4D733E6604A003C804BD380D6046469E310AB9B07CFBB605A32DF6E1B15734F8C2580D792AE5AD45C13C37D90D893218FB7BC6A449161C0B91B2FE8197C81929EC8823942A2EA8F7C04A307249CD3295B6B529CC87041B6866E9F358B5EF30486D7CE9BB297FE73B2A0BF7FE5D4F7C56281DFF8CA46B5F1DA6A14A15EBE6F6D7DFC4327834E655CE52C310B6DD6D72A9D948A930A11FAA6E57A08A6FB873341A3F1211D0396884C07F785BF4531839AA77EEE2D5BD8D1B767602C01F6CA35FDB0F6A3967C367F88762FFF45A67A4E75C16F744B6E6FBECEDB03B346EBB18B1A35D0F2CF387277CE01F8068DC250E19F0E37FE36783C0D4FF4A1292577DE8F3E81CD769B2D22EAE286E75756ECF31E56B00A57DB2C17750909ED9959946C86E25112ACFAC5F526A331B5E49DECEDAF38EEFD5D5368A8539E49A0766C22CF5F713E6EE058E9BE157805A521FECC934987809B9C5190EBD0E709D1B2EBDB06F925F3203131171ABFE76684849C0A82EC8D66ACD60A24794BD39C18782506BC7F9F7DC6B1BC7EB2D70A3FD7AEF3DB81568C5F6513161D8DCF0B9383DD97207C186572449F7B55806FB564723729394C85291E01C5EC803D8FD2D702BD9F84BAC47E6E659A3FD90D04B4F53A01DEF302898D4EC430BEB2936C70B976355DC2A68D798EDE02F534872E369582E8B4DF771AA3FB15C2602F2487A21EE9DCA0C2ABA12ECBAB2C8B49939180C3E305336EACFDC339F502EC730B55E0FE4227415EDD151811D018FB34839DCDB684C9C8453F681916316DADB8BBB025A6B66DB0C6315C73D0654113CE37FAE29DA59A893C4C7F001DE15F0AE4B59C211EE59808021DC7CCFC2BC8B2C15214B783FC55E8C50A19ABEEC8093D82C3E12058B7023AE561384D9B28307EC60D004BE81512B0D03F02388FCC2878832C1F881251BBD73D3245336E12653445B6CD704A796A284A7A7F1F7F37DD9D22C2B2BE0D3C497E2F25CB95933D154199A32D4971965BE442C914ED7C42F28D33BBB61684AC719EA5F4D7FF7202E3D476519B3CA236A143B1DD22B34F479C0519531BBFF5E1E1D8330B231D588AEFB2BABEE0A1BED4A1D775C5BD5177A8CFDAF83E5B4CE662418D4A13FE34D3875E9EA15BAA45033CFD746673AB16FDE39F31BEF02051CFF7DC335C6B9DD8CBD17CA9B652F01AF2E3044FC3B1F15378A967F023DAB2AFC2CFA577B82DA875E1FAB014728BD7A8948859EE9619EE02DFC85859D28DAD6B8B2AA72F7973D6709D1DCB0C625084771F3EAA12D4B6D091E6E5026845F0C30FEED6BBACD4A9B5D623CA247CD6622D1E18590E5EF3FE9A094263E886E567BD1AFE24D7E263C5B2CDCF03D1FFE2DE85D7C81A7634066B30E0FF49B71234DB9441017954CB05B8BB72C11710A55041C737AD29A58B9EC6E2CD871B56976C389133F45EA4A6C39545AD15BAFD9863A333637F7AAD613BB82E61652A00BF90DB3FA1B4205198A42151DE6A3500F0A770AF589AB63C01299A28F94B9395D652866BDE7505BAD85DBB2B9D56E43D02F679F94B4F0DCDCAEC1487E18B89F96BA1F1890BCEA47E60FB0165092BA684F8381625F83C86FA90F006";
    keygen_kats[2].expected_SK = "9C17C88109B6927D423D887BC2FC24A5C4405C8E736C1C9D9A799C5CC09DAC3B0AC8866103C621D3464AF8A7E67C30C8FA7F66580CDABDB9E6848E611578D0E85F99D936F0B17CDDAD87C4107D0642F26EABDDE9732CE11AE78FACD7532C2868A1A29A6B5A0CDD35F4EA2F536DEB14A7146F4E94F723B69B976F4688FE8B5D22A0B281D1426D18144D1A066403A98808390E010241D32428233764A3C220190322C8C0405A9265C8B82813B789C9089211082AE4B464D018300031644A928812A52DC2280108C58559A86111270912080D4B384621B144994268C0062999228D01A511A2C46882928C24B70D81168ECA0465D920289442329CA00924356059348EC4C46D23C52123A425CA10921441240B424E02C94C6094318C082908260440046249304A21154002180DD282294CB051211406DB2480DA08012125661B96641819125B9649C9406C180004090380CA1210D0444EC2A271D822694B2091DB8251E0A00D0C9788D044091BB020C3C04024C7251849450AC84001164D1BA96960A691C2B2288284818BB44404B90C9C4206D8063198926098846589240800098209B349A0286CA3C428C1145198222919266109A208081152E082895CC06423A641C408721126321431122231700B15868A16426480311B156E023702DB4491A130804114200A119098142519A1519814264B422C0A878DD9386402B33080B25104B785D2120D11C44864A88DE2868D1C2090CA940D0C15500A188011870513988D94A265CB164D1486418B168C88002D14C680A39069989431514866C44286A304302449048C962C0312806124456312806182098B300699A65002942D08C44124C96C000546C2B6098C0025531872CC108C13A0458482080A972554C2886342859C3049CC18929AA82013220AC0282694367049A60850C850A0B22C60B220A4388D1A128008346190366C0094700A0912C8302C41B66859B669D4C2814226699A2404542442A3245203115123234801B2001AB24843B0615806890AB66811B5641230841AB88DDB280A2437645A262164340508075200B7689B988DCA164810B9440B8490E0A41011880494184013B500440060181469540050030864C40062512030C42200C9828900496CDC96404126051B87245036495006029116449A105213A62C528224214690D4364D24014044B628D8264AD0A26C82288AD4C66920A36C49A40440068E63B405141168E0264008884419158C19C62994966110868041C43108458949B030A102851990041A166A8AB631C33085DA1672E2028E119711E128810C8388D21200CA164419C52544468D1134615C946DC0485154808C9C045153040E09380D110248D814880B88719CC60C64142812854801938DD894890284258312698BA828C2A690D4264504B57120468D21462E410241A3C0082030028B442C02264849024D530065CA24465904460A290E11A460D0A020D1140D130185D4B829494684989081DB2290D9B011C4460209182C63484E4314001CA24450B20CE0C48C09C98C8AA28011B06058C20914B9208C384CA0A49124271223112C63807102B31048866DE0882D03488C61A4895C241143282541409118286D54261191B82CD82069A4A229E4304153A20D08C1400182694A440948222D6304066434212490648006418AA40DD094690043819216649408486094715CA24D61248018B8814194200AC650E1468A4CA65192822844140D4B2006CCC84D1C3460D04069208641C4C66DDA904880A2111BB44CC4926DA1B0080C11724C204C93406111494258948920388C89982504A68813412699B6458C148060288A032402A442658AA82C1AC5412288705C882114A78C0A447241402C88180012B48C4BA8640A934CE184400A984DE13070E08404230900CA326249846400378492B08141A629C20621DB162409B74DD9A28D1A8208A3388483B60C8A824D20B48C4BC82C8100640BC4850A054E84B04CC1204C503851131305CBA210040002CCB660DAA8084AA091121121612401D016920CC950849804DC803081A465C986301803321BA1681AC904D9062C042149CB480EA11088D00802E01086D9346C22850C9B420A122948DB0089CB3088D9940891343294C8051B940420226010849114A58CD9341101355020C361A31682630231CC3881DBA809149349038948134210A304094A2688956D861BEC7549AE8CB7B5AACD88780F7B1D1597FA1BE27973CE28C4C0E9F35194AD0E2DF62E622B75E06E7E21AF5FDF3E4908FBA7D0B657FCE0A512FBF13D3C83F16CD3BE385BA075CEE26E68A28502C3C097539430E8F19916B44E53AA7742910B719CF4969D5EE2D246F5CA207AEFEB037E7CCD592094DDB72621C5937813A5B324ED4544200460F4EA7744DECC6D182A604C142D6212EB6F9F90B1AEA0F89EC07D9C083EBE1FD78D3C4C2282E1D5BA47064E8DFE71ED9A7FD7C0F95481F3CF0610CEA3FAD5C4E73789C70AF963A1DFA6DA9DF610BB98630EB4419399AFD1412E0693E33BD24381050FF62883D65150AB1DD0C67F443E5FD247412DB729D2E58453C770F934C475B89B458111DC6268F1CA0E9D143E7F0570D22AB5B7BD9446BFC7DEA9F06383FE1A0BD9E644CAF2B91AC44BFD37DEDAB4237990A3AD448715940001EA30E7219172B64D86E85C1FCA8DFA922B61819BB4BB68FFD44970FFD9CBD6BD2F09FB12E5265A5B0F919F6D4D6D06534FFE792CDF6882DA5D4557B51AAAF3A80A8CEA69E8678E66D1F47592BFF128EAAEBF38C70E8FF7AD31035DA28AF239FE245D2FDD4F853029A65399D5E6B6F4F4CA2D862B62AAEC8EFCC4B05DDCB351DFAAF1F7E7ADD9AF9FF44D2E2A384368200217F48DA0DF5013BECD2462D4BED2359FE44D9612EC6505A76071E116AB5F0F1DE88288DBE97A8B0EA32B9A6FC53695972A8F6B33542457C30C553DE91B118B15A6DB2D3F56FB0CCA91DF79741AF737E88A88A69424F7192EAFB981DF8256989189D75E0C7183E3ADA99CED3913ED35DF5AB82C8FD07D7B67DAB7EF443DF51D82FE87F8CAE103713F88E9B73F649B1D3C8589B71F06517B18502CB230EC27150C072D985A98790DBE1F83BD59421D19CC9E23D845C50CEA8515690944950809CF95FA636AB3509AFA1A7ACD2F6C346CD76362D15907764749F3E16C8BC84186E1FC9FA120F49859F7E4E6C75F7CE19C9C129C72A7CA129D10AD8EB9650DDB304F5F02FD7257DD8D71B97BD9ED47B9111236E3B706AE4800401B77E1E5A541E44DC1D686234884A5F910AAF16C8D23E593A307DA8F1180095D7A707566E9CBB125751499D748A7E1A78108B93DCFC165D2906A1DD9AAE8C5BCFCFD1D5879A8E30B6FC3EE38F470428E8455162261E7FB6F8D5BE329C0FD494492C296DC8A78128478F88BD6E1B2CBBD731ADB947300A82DE410B27C87180032AFBADEFF276BFDC0072179E36053A3F4C031FC2F94116938EF7B2A02CDED2C4C101AC0CBF0F0404BF9246F1E4B71EE2EA0569BA6478C4929DE40C56B075432203D8CD2C0EFAE663001CCB0947CA073C0301A3896793F7FDD0248F7CB4CDB184408FFA24AC8016716A7C40572731CC95DF6954A94BD2E507FCF71A8E250124E29313ACD6AED2EBBCB36ED59F102F706D5E1B79DC3D956F46997B4172C7FE20F550CFA0F1508312CAD73AAE7AC30BADFDE7D2A8B2ACEEA2FC564354276AB61A8F2D6A3CE5D43A5E6496894B66E72DA30370692421D267F04430397C3B9293F7EB11C107C2D2BB007EAB932BF25CA65D050CD061D3653BC1B25B5AFDAD7A9EA9352718CB9584615D8670CC61D7C165D778EB2766930470AC115F488C3767A6B80D987EBEA29839642720275E20602ADD280FFEF51005BE2AFFA3F69BCDC69C7C40FBDB9F8AB2C57E8745A9CA2124FFC3E088B5564C088B71847A2AA574A4251C1F5ED3F02E22A85BFB1AD2B137477439D4BAA4DAB63644A44C0CB121478A2D91E2B7B9D6CD02968EEADCB51BC5450ACAAA81EF9C1A05B475DF46C4D6603C371D6AE3A1E777A789E7205EF7AC574753F60493B81F8E0AD527A6A561F5C1723EB7E9AC1D82658C00F1CC538DD8E5552366FC9A34D0EEE1EEB9C4228C58D2D7132E3599686930BE56B9A59097B2238AC49FF4F6A9F893FBA76F511C6A6126686C0BB6CB946B0D3CF7DAFAC886BEC911564332E773C10ADFFAD490B94EC6545DF90CD12695E79936A7CE77E66C3F2781F6606874BD2E1379A8610B0BEEEF465334A455DC2887D8B35066B496856A5500AE079178EDD320A7AD2F0D350B0B3E78EA658787AD5F4CDD224340E93A06996904F9D5EA21219B871E21DD3BF7BD3BAD750048702059C86584B0E8B4EFB144503609D021C1DBD98F04C84BCE4304C834BB502CBA56A6AAFEAE643F76FBE439033D13F5FC93D8D852710C3CCA4E2507CAE51BB8779C622AE8197CAB5E51C9D11BD38BE4145CE12BFDA8F8B9ADAD8D8033D38143C92ACA69D5F72ADACB8D6BD10D427726D0F51AB7114A174E5187B8F9D114C2F4FB768EA80F74A49CCC642F5DBB7CEF2DAC669E250451CB9AD8EB2A7631E6884934E2A25FD710F3E47726D7709BC89800C6376158917026C299CDF76976624AB877136A19ECEBBBC1C36DE60EBB3CCBD43508EE6CCA750960543C16A0EA3676CAD076DC3464517FBB3B2D929AB2FA80FC0B31BF2026E4FFDBD2C20D2DBB8FA09BD88CB4B3CC124CE260BEDA345EE0232B2034AAE1E1918365878D4A0BA98CD4D7011014FF7569CDE130389A7D59E860AEF59BEB4F4D3259C1B092E68FF8AF679327F4181F6476D54D933B7EA376B1D4C0564D204CBE631C4AD3DB45F3A7CB894AB139BDEEFBAFB6EDDEF0DF6F7FD5EF140882E21CE59AC45417686DF7CA38AC90A7B44DDBE0F085CC397B3B65E6D2524CB2A6D4AE4BC69911CFE84465C9D6B697D28D84C8C28EF60ED5BC34B0EABDAE529CFF3C00F0C706584C48B565CC060A80F6DDB0DAD0799B8907E94B0C29A4E7A8D6CF0C5750DA5EB717B30341352E6046420C7A226A1935BB7F0D25E4067E30B527A55BF410B4335063ABC9BC76A5D885882AF728AD934BC7E55553B9ECA69D97311EB3CFB1DBC28891D3DBD954084E911DCBEEC1056C502385C8EDA9B4ABB93E623132084C5950FCD44725BDB70C9B9187A30DF477E128F143D870A7F02E5D2F20A3F1B034FA05475F58D98A6D8C22FFC0ED3792A1A2DDF00F62CC03CA04060BCA60EBB9CC27C2BB6636BBA116CFD03BB196D85DEEFFE0C2D6359129FE1877F723EA225FEB1E995A34B9A3A75D1E6C0786590E159CDD62B39D084AA5BD2EBC4456E694054922D4FBCBD5335F7F8448ACA08E650D296D45F3511365B5304F1359EEC32E4616C166F938F2F36C790BD577402C4A605149A4B4F8E1A101E97E22AEACFA89273B3C1824B42B0019AFE8C4ED8B7F6A265573E11AF026464BFB2C78532C0AC303EB5D36D88CC33F528E56310300D52481BBB27B7F8C523DC036B2D1A36C002B98BF5F58B4254D097DF7912D4189287A14D7AC1A30691BCB53FB9E86056852075B7278E4A50F76EBABC11761BFC5D2A86B5995B1CAAFCCE5F5B3BA2C195B692743B637E424AD4072C4B5DC6BE4A3DE4E041E72C64FFB9AF9C66353C5BB2A3967830B9CFC9AE5C632A14BB32797BCEC4A595D8761524026F13D237B165CA4240D4972287ABE72AC7F419F37E99047F17D5D9DB57C508AA0730D6D9D2049E19B1EB3C7EFEF2EE719047A777FD281A0960C09BD79443C5891AD8BCB1ED643B9A9F1E66FB5C7EC6DB926CD73DDFF4D39B15E386AD92170C4F678A7BD7FD6EFD600FE082A64AD91E2EDC675DF911B531074660096E85C66005318A3B85CF7E1C5D269C5BAE4096C9E05145C01C9A6294A50B3D4707A93254B0CDAFAB7B0ED1CA6CCB3DDC1FAA5304055C41095C503DD79F86A499F292C473C3B975DBBE53216C85D42E3E5A819E1A947639131CA18CA7831091D64FECA2713B8BA5577BB6B7FFAB6D376856A4D38856651EBF90929784436EE1F09EC9C99A2BE601294AC1C7ADBBC0EB050BC3F728D5D0F3D4831BA4DEE0E4674EBA6C2D26944029B8BBF90891C37A69DE342EC829625544A82C3FD8F61DBC40ECCC6527E06C26868B33BA362FE4E85FD8F76132E9065F6FA1DE7FC0CBB92A3306534AE9FA01256B24ECC2C63854D3F46284D0EFFEE19CE5B7998DD8DCEB38FEFEF074EF35A3748A9E44AB4F75F656FD08866DDC4F58252B25A0232180E8DB2CE8D346A558B03DD71B19D81E5B23BA688099DDAE1D10BF52932FD2EBD360E653BD4C3A254FA4B71F2859757FB024B14356BC00DD2877AF29BB57ACD812C22119F8CB62BA81C946C36B0D4CBE3A1B4810FFB27A47096108AAD74A5A0413D2A1B85286569853AC230BE9E34C78C84FE0F6269685878AA1246A55F37842584EE302301941B9A6CFB8BB4ABFBF3DAE55AD8ABF6CD6CD7B2C881DF7D5DC264A5F61584A990A8D1CCCE1C0CC05881B4358494283964EEFA16E9A47586FB9ECE3B39777DC6C1DE6931C5448C0AE2D6C51924D7F6BFBCBAF485F0F22FA2228A162C13240EB64C050F2EC800E937FA97C77E2854693A4CC83E1773EBA74CAD800F4AC6CE461C9693005BE0B3C288EF1898900466318B96AD247139E5E8D8CCCAEDD20719275E102F50F1CA019692642092CBCB21210EAE0DB708D96E50FF249E6918A628B7834BE30349EDBA515A46B0229E6E7AB1A88C25A7F6A3BDFA84EAAFCB52AA1A143FB09DF7CBF6E39FE1B813AD64FA786155C298D9483C2F9B39CF46F936AF6B95E3BA82356D7C99EDEE47CA00C3DF9A80E8DE0F246C5DE4FEB6C55B457A59CD82AFF7A60E3100D409E3EEBF2E695DD3D047CE2B35D3820AA8D4D7692C299C00B78EE7BA40DE61560CDE3FA77BE3AE68E";

    // Iterate through KATs and validate
    foreach (keygen_kats[i]) begin
      parse_hex_to_array(keygen_kats[i].SEED, kat_SEED);
      parse_hex_to_array(keygen_kats[i].expected_PK, PK);
      parse_hex_to_array(keygen_kats[i].expected_SK, SK);

      `uvm_info("KAT", $sformatf("Running KeyGen KAT %0d", i), UVM_LOW);

      // Wait for ready flag in MLDSA_STATUS
      ready = 0;
      while (!ready) begin
        reg_model.MLDSA_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", "Failed to read MLDSA_STATUS");
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("MLDSA_STATUS: %h", data), UVM_HIGH);
        end
        ready = data[0];
      end

      // Write SEED to MLDSA_SEED registers
      foreach (reg_model.MLDSA_SEED[j]) begin
        reg_model.MLDSA_SEED[j].write(status, kat_SEED[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLDSA_SEED[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLDSA_SEED[%0d]: %h", j, kat_SEED[j]), UVM_LOW);
        end
      end

      // Trigger KeyGen operation
      data = 'h00000001; // KeyGen command
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE_FAIL", "Failed to write MLDSA_CTRL to trigger KeyGen");
      end else begin
        `uvm_info("REG_WRITE_PASS", "Successfully wrote MLDSA_CTRL to trigger KeyGen", UVM_LOW);
      end

      // Wait for ready flag in MLDSA_STATUS
      valid =0;
      while(!valid) begin
        reg_model.MLDSA_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLDSA_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLDSA_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end

      // Read and validate PK
      for (int j = 0; j < reg_model.MLDSA_PUBKEY.m_mem.get_size(); j++) begin
        reg_model.MLDSA_PUBKEY.m_mem.read(status, j, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", $sformatf("Failed to read MLDSA_PUBKEY[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("Successfully read MLDSA_PUBKEY[%0d]: %h", j, data), UVM_LOW);
        end

        if (data !== PK[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("PK mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, PK[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("PK match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end

      // Read and validate SK
      for (int j = 0; j < reg_model.MLDSA_PRIVKEY_OUT.m_mem.get_size(); j++) begin
        reg_model.MLDSA_PRIVKEY_OUT.m_mem.read(status, j, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", $sformatf("Failed to read MLDSA_PRIVKEY_OUT[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("Successfully read MLDSA_PRIVKEY_OUT[%0d]: %h", j, data), UVM_LOW);
        end

        if (data !== SK[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("SK mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, SK[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("SK match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end
      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end


    `uvm_info("KAT", $sformatf("KeyGen KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



