//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef struct {
  string ek;          // Input EK
  string dk;          // Input DK
  string msg;         // MSG
  string ciphertext;  // Ciphertext
  string shared_key;  // Shared Key
} mlkem_decaps_kat_t;

class ML_KEM_decaps_KATs_sequence extends mldsa_bench_sequence_base;

  `uvm_object_utils(ML_KEM_decaps_KATs_sequence);

    
    // KAT arrays
  mlkem_decaps_kat_t decaps_kats[];
  bit [31:0] kat_ek [];
  bit [31:0] kat_dk [];
  bit [31:0] kat_msg [];
  bit [31:0] kat_ciphertext [];
  bit [31:0] kat_shared_key [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    decaps_kats = new[1];
    kat_ek = new[392];
    kat_dk = new[792];
    kat_msg = new[8];
    kat_ciphertext = new[392];
    kat_shared_key = new[8];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // Decaps KATs
    decaps_kats[0].ek = "39690870B765DDF5A0B7092773EC1911637E8A80307A865A24E3012FBACC0FD431D12A44B38CC685335C858714026187E8F641933291CBE0B678D78944B17D7DA605DEC011B8681E113701C0074553156EE11530A4B63B8FE886637B524DE2733D039591230CD90C1EBAB61E3A5762E46B4E6067C6C4B280F371A3D8BB6839242DD3E381B41A3624396C2C557D1809934A901D8091731A43A32DA32EC9FA860FFC4AD09022B944C654980D2F928773B5BBBE048A21DB3F67167EA7F2B156246014ACCDC24455F5D1B0F7171D29CAA43DEB1CE32513078B495AC09C9B6793497BB593570CF8AA2D1F7549E5D54FA5A339B4281C90D75A9D0186B7322129B90B1DF6A39892C60A613D55E4A46EC07B69B6AF96255617C77951958A15B71DC48075562A236AA325008909CF75993CD58AA81658750985FA593EF6C0400BA07BF119C7380B1D61751A4390A398B6205A6895A857A463EC931FC262D89B069D6CB3AC9BB4E5272F35CA612D8346B65427708186C9422A37332B9955BFBA7080454CB5972397839B5465219EC6024D08A46EC4B29A15249653F413FDA1C99E82C144E7BCD9E17C19C2C3D43C4792F91EA4D8487567392AF43A513480975959E50CCA55DC89AB0A19A313B1B7E6ADBD7A1477281BD128B2C0F867CCD13877248E5844882F48B878E536D5208716F11B75051033E9A30DE9AFBBA66305E1BA265686B29C3186FB3CA1952936FABD2EA931E0D74E4D849CB685BFFC38C9E29559DE6AAF2EB4017C543EB9D59732B421C3A5CB5781BB60F1A953F07D7937B3651305E1D46E15569321721E310494C2EC16C843B3B4D9831809065BDA8F4E5A17E80123312C065C03ACE623AF5589CE361C913BDA355A031E42C54EABA24AF3F6848E6C4932427AE2A09D25808BDF0288D4C245EA2973C261CB29A6AFB13C6058A3A19F11673A198F86A251113837CDA27F2304A1E3D75C8BB88E6C67A006CC63DAC90017B865DC0268EFC53E2CB75CC6F1008B34839CC80B26A019440C0D34132BC4690519131DE15434B730B3A2492F6EF6471CF1C5568463A3387102135EB1A8635F0A63E33176914B40CC2494002C0E19C38A0D97C0CA5632261519193030F33ACEC68125D33C5AF26A9F97B1B181A00E4E9144A2D4811D7654F9B958CCE126E030A7FEC045A0BCB82ED40509643F3F5736B652116A4008EDA65FA1895EC82390C2713B4303BB6E7B4B416429D8ABBC497B98907224D065B3DC5A017907BBF7079E08B770AFD059A31A30933580EF49B5C48B0ACE675697D6B1041992DB62246092376954980AA03DCFCB5ADEA36B0B2138AE349D5E270F0D83640BE9885CC9371C6490C1F39959C9A192E584DFF9CB2D8C2297B117B9D7627AC5B2D29335558718A5A7C34564B0C0A1105F0A00E0084ACA185C5A54741E4B4053A431713678F5951D3FE47E0719A082017AB73B892EF3C77ECB170BF386AB36C89876BC8AE67B0CB82EE42793D9D7435172043E8CA3A8E1A83197891121932A0AB2EF46789EAB0BEDF5A5707A4B10035BD331B01E298370E112443A48D96CA9503832E3495DD2E571374C1F57B6B9A0A074AA29736C488FE1D823662ABD3A379CA43007DE317392D332A6826ACE381AF4C82C31F7C781788C705C4E6F06B1488850AAE55B6872731570444DB49AC9A53E9635816C1C537D2430F922124317592B36A68685859EF334B2782A5072A661C55C39294975572319474DB4E33DFFDC5E88ABA83B6B8D468753C88BA898DB116CF0415DB41C17D346462BBAC4A44207D0C93A4B71C8D00D47B969C690ABB371C0BBE1A367A3046643C466C867E341805EB435F8316358F69E6A4976BB54ABD90AA963B52BDFC93BA27C833BF5CCB4A2CA5BABA12D70016ACB875582416BA1A82246CAE8489647B36990F9128E350407CB614C926E492BB6D78021E73CB54641317FF282B9436462183B9375A5D32879355A96215B31ACE09C93779240260EB8B974FE049407229B808B7818142C3A071CC5561F56593E7605346C63817FEB0B836ABB786077BC7A7E3511275C160BA9017C57774E9503048C29B959F5C9E354A8E137CD72C873AD1978F69324DC282504E0A221FB1B740004A63AA7A2D33E00BD0DA29962B8F30233C78317F22CE7D068F16C1722994225E800491E05723201D81BE63E10D05502E1FF54580492D7DC5682EBF09E85773B4E61";
    decaps_kats[0].dk = "042C24A9415FEDEB4932F34EC4D30562112740E60221697FFECB24DA0888D71456CD7924E9669DB01511EBC3ABF6EC2C291146FDC90ECCC3A270BCA938332D1A09019CECC35F8C7F8FC419622185D5B734865C2DD4A634D081B098EA311A029169C973B643C062CC7E31D73876731DACF830955A7F73B9BCC9D6B6AC4168F747885D3A3C01CA4AEFA20EF5B55FB176AE90939C12002BA9324752AA2A1DF78F3A6834FEE50B5165A4AE0BCAAC06BCC6A99E94A69E81E65207F52AC11088ECBA901612CE8BA67788CBB69D137479F3A7FF2513FB8320CA946DDCA952D63A67A5A0AB295249C76169A5E09915BB7DFBF2C876C897463C2B9A973E5906C410D7A04FAA0D2813C48CC5BBF733C4A706139A1990FA9B1E78A98658364250837B34F8120746624AD67C2FD8C5D92C3A0FF300C094988CB077FA65547E55940357AFF18266CDF511E74069E4A85797564800D377ACE053FEA919BBC64869355F0618813E603C1E5B552D624D37924D64B83471C6186EF763E9F319CA41009133360D45CCFB3C8667D3ABF1EA7CE4393683EC9EBF88B3CD3C3D30A6BF66D831FE235CB7E95AE14321FDB76EA59345DDC21D4F6C5D7F5105A67C9CDD6818F07223EE97518FA666E526A0F489677B004705770E5F2B68AED90A1E69C54BD0A6901C766B3477C1DA346C95217F5B8A4475B2D6C0A7B2708A4F519EECD1A67B6A3765003C1EFA308479ACB7584B4D389AA0F3200578C2836AB4AB532686793BA9C078A1EC587755C6DFD5B7EDF41684A3465CAB3D0DE80E7B83C16E7953C7BC7A313B2DBB68B204EC7669730AB3ECAF610C9158230323A86A4B8AB0172A8F7E92825F8C7F1362CB4CA4A4ED1973C1D620120A638EF88EAE78C11F90B0560809591293A3DB5D5409CE3C38817D1C917EAB8050E8C69AA6C8F33178B01A9E6CD31DB60B15FB7445A4149264D984FB86AA5EB6A77F700E7F5890E1ABC2C715A45B23192BD2794ADA65BE8835F2DB9563B32D64B65957224DCE30726A6368AF7A3E016B7712A4671DF346173411EF93119B071AA19767C64474DD317174C1047CE60155967982E661BE441C9363A1CFC33C7CA7CE6A620CB13879D75C92E322C50C9C0C6A041492EB5ADA1B267FA0138B63A3EFD8A2C3F9330CE805F5516065230E2B9C89A2AC3BB0C231F0F8A55265CD143C22DB873FA90068027A3E21275431922FEC6AA8E5F544A3389F8CDB051EB849C5250D27D63D8F398DC2A172E8016FADB223D47B9DD55BC01230400995B3CFA51B16C903EB8B4E4A9704E748006CD1710925B75000CCD5724F3CD81BC68C9364E36BFC972842274DFAAA2D85816298C51B656092522C895B9B1B19399A1FB28B4534952D51C6EB16CE12A16838C64EBE942C90A06890C3246C1800C0F5633834932744B8B5478364D7272F80C97D5A0E19A37E6B182812A0604B5C353274A139DA2948397ED14286F902B5429B7FF5F4C84ABB3FA7E1A805974C89AA07C906109A73C7B1B0582967A2FFF137B289CA0AFA3B07C221750A7CC960B6A679B66AA37373585F8459A7E3725BC718382FA03BD433AFAC481BE5A09B6D2075DBBC9C4CBB92BC915090D503A5ACCAFCC2A360142765FA2599A55DC05A6A2D5300F863BFE7DB0574A102D76C1773A095F3828BEAB7B0B945B19D0C288294B6ECFA551FBA26FB58BA8FF39499ABAC74B990995592CCE5A2EC8625BCE26C4360875B65C1D1831A1854303CE780198551015C2C62F9AAFB70B1A15834D467A642B180BF99393B22774E0B3706421A7AE2CF41281BAE15891E429F74314BA63B02E0A661C2891EA947B7571CC47ED749D70B0595203DD7574AFDD6AEDF8CBE55FA5D495362DD534C37B926EBDA468A48CB701C0565A81994C4AFC599223AC963677C9663211D7B8698D533673E8356C4BB6F77B6CAD027395270625F0A80D5B5A881E61C9553C165F9CA2B309BA7B21CB516392955617F9884A75BC797F1098D226F821985077669753018841A9F290170252771D14BA8FB5BCDFB33AAA17B6032D3540A08B85846212AB0C40430A209A7244420B5A81357FF669A4944291AEBB50ECC3EA8962236D2C4F8CC0354074827D0A37EBCA11292A9D41A7F06D97C37C2541593AF33AB431935CB4522370651A784CC5529CCCA9296518BF87239690870B765DDF5A0B7092773EC1911637E8A80307A865A24E3012FBACC0FD431D12A44B38CC685335C858714026187E8F641933291CBE0B678D78944B17D7DA605DEC011B8681E113701C0074553156EE11530A4B63B8FE886637B524DE2733D039591230CD90C1EBAB61E3A5762E46B4E6067C6C4B280F371A3D8BB6839242DD3E381B41A3624396C2C557D1809934A901D8091731A43A32DA32EC9FA860FFC4AD09022B944C654980D2F928773B5BBBE048A21DB3F67167EA7F2B156246014ACCDC24455F5D1B0F7171D29CAA43DEB1CE32513078B495AC09C9B6793497BB593570CF8AA2D1F7549E5D54FA5A339B4281C90D75A9D0186B7322129B90B1DF6A39892C60A613D55E4A46EC07B69B6AF96255617C77951958A15B71DC48075562A236AA325008909CF75993CD58AA81658750985FA593EF6C0400BA07BF119C7380B1D61751A4390A398B6205A6895A857A463EC931FC262D89B069D6CB3AC9BB4E5272F35CA612D8346B65427708186C9422A37332B9955BFBA7080454CB5972397839B5465219EC6024D08A46EC4B29A15249653F413FDA1C99E82C144E7BCD9E17C19C2C3D43C4792F91EA4D8487567392AF43A513480975959E50CCA55DC89AB0A19A313B1B7E6ADBD7A1477281BD128B2C0F867CCD13877248E5844882F48B878E536D5208716F11B75051033E9A30DE9AFBBA66305E1BA265686B29C3186FB3CA1952936FABD2EA931E0D74E4D849CB685BFFC38C9E29559DE6AAF2EB4017C543EB9D59732B421C3A5CB5781BB60F1A953F07D7937B3651305E1D46E15569321721E310494C2EC16C843B3B4D9831809065BDA8F4E5A17E80123312C065C03ACE623AF5589CE361C913BDA355A031E42C54EABA24AF3F6848E6C4932427AE2A09D25808BDF0288D4C245EA2973C261CB29A6AFB13C6058A3A19F11673A198F86A251113837CDA27F2304A1E3D75C8BB88E6C67A006CC63DAC90017B865DC0268EFC53E2CB75CC6F1008B34839CC80B26A019440C0D34132BC4690519131DE15434B730B3A2492F6EF6471CF1C5568463A3387102135EB1A8635F0A63E33176914B40CC2494002C0E19C38A0D97C0CA5632261519193030F33ACEC68125D33C5AF26A9F97B1B181A00E4E9144A2D4811D7654F9B958CCE126E030A7FEC045A0BCB82ED40509643F3F5736B652116A4008EDA65FA1895EC82390C2713B4303BB6E7B4B416429D8ABBC497B98907224D065B3DC5A017907BBF7079E08B770AFD059A31A30933580EF49B5C48B0ACE675697D6B1041992DB62246092376954980AA03DCFCB5ADEA36B0B2138AE349D5E270F0D83640BE9885CC9371C6490C1F39959C9A192E584DFF9CB2D8C2297B117B9D7627AC5B2D29335558718A5A7C34564B0C0A1105F0A00E0084ACA185C5A54741E4B4053A431713678F5951D3FE47E0719A082017AB73B892EF3C77ECB170BF386AB36C89876BC8AE67B0CB82EE42793D9D7435172043E8CA3A8E1A83197891121932A0AB2EF46789EAB0BEDF5A5707A4B10035BD331B01E298370E112443A48D96CA9503832E3495DD2E571374C1F57B6B9A0A074AA29736C488FE1D823662ABD3A379CA43007DE317392D332A6826ACE381AF4C82C31F7C781788C705C4E6F06B1488850AAE55B6872731570444DB49AC9A53E9635816C1C537D2430F922124317592B36A68685859EF334B2782A5072A661C55C39294975572319474DB4E33DFFDC5E88ABA83B6B8D468753C88BA898DB116CF0415DB41C17D346462BBAC4A44207D0C93A4B71C8D00D47B969C690ABB371C0BBE1A367A3046643C466C867E341805EB435F8316358F69E6A4976BB54ABD90AA963B52BDFC93BA27C833BF5CCB4A2CA5BABA12D70016ACB875582416BA1A82246CAE8489647B36990F9128E350407CB614C926E492BB6D78021E73CB54641317FF282B9436462183B9375A5D32879355A96215B31ACE09C93779240260EB8B974FE049407229B808B7818142C3A071CC5561F56593E7605346C63817FEB0B836ABB786077BC7A7E3511275C160BA9017C57774E9503048C29B959F5C9E354A8E137CD72C873AD1978F69324DC282504E0A221FB1B740004A63AA7A2D33E00BD0DA29962B8F30233C78317F22CE7D068F16C1722994225E800491E05723201D81BE63E10D05502E1FF54580492D7DC5682EBF09E85773B4E61D4ED29FB6EEFC6279C24822EBB0FE9B69246931ED0467352B7E69E79F47CF6EAF36E9099A67947E97C78ADE6C5B36316336C025F16E7335BD81A3158D5AFC87E";
    decaps_kats[0].ciphertext = "FB25DBAFA2CD7DCE979BE90E31179FCCC24AED8A86D60C3B84DD6F701B249AFBEAEE926F05859F818CB356FAD2593B6340B6E59480D7E78E54C54D3178BDE122F0D3010BA5BF2B65468220088DF430E1974416E12BF5B3B3EACC2A3ABFC038460D83257A8CC7F4283C6B3D0070DA8C8BCEEB976C0D708D056F04C86E35B81E99162AC72618F3A39832FB90B378DC914E0732F3140049B149292C8D00ADDD9C0522F3BB1775074AAB4F1E279B5946E88D7C46CCFF453B55621817B8411E24BD0B90BDC275822A8164BA11F9477AE9B03DE7DEA010100B164E02A91F0A27B84B585CC48D4AB84B0A1727454BBE84B1E8B723C2BC7A4EFBFA657F08E7AD2670CDC497D534F307246265C89AB4066E2E1101282A328E00CD1B58E4D23F24CC364CD92F891F4815FFD974ED36C4D29E3C0C7F302F0E912E1080222134ED6C973C8635062F63A39762EC96C883A012F369566B62FA5AFC142E1E284675E7C1EB4744533EEC5DE95AB8ADACE27259DDF76553B482CDB83F1414C66307389F82A51B949AFACACF5E38D677456A8CA1806CC82E3BEA884EDC7B4C5ED66007B143F1A19AFE1A5540FA69F999FE86386FE1E83FC0E57423DF35E82749ACC856D3F05EFB959169CF03C9CB3D11D88FBA1F85979F213FC59F084B01F4FEBD9CB560C0F969F8F021C30644FC8721CD12E2E2BB0014B39D9FB4916FD38C6F8D9B02D67DCDA44332DC519528A86DD5161E8B4C100CDFCC58E3E05763E9FE5E69CC5D5C28E6D2AB24A4BF853264A3CBDAE0A72AA380D37CD0D306770D711BBA1D55A13EE7CA01702556B57BE5F002FDB6CE00DE00CEF2869092803CE44F4944A60CCA2B30978F39FA644A96A66156705EF1E473BF38EAB139AEC783230472CA49D071A817375191B891A9BF63723BF02830D1F443660B33C5EBCEBD8FE04BE4812409E82AD48A21C50C241CEED5126AB40148ADE08E12B381623E5471D173E2722DAAB9085915026088537EEAD054C7207FFA1B68F9CC75DC34D540B7933F78FCFE5728841AF808C0FB9D83F6A80EBCE6B51534370DB55E274B74D216C249759F80D9494EA1FE0AD058F057FE3C72759F5F787B35B13C3FBEC4B730244C0056FE694D801C021DFC1F179FF6BB8435878EAB8936FFDCAD68FFBCBEADD1BACD3A6922759DA01E72AD933F34D10F29D74470F70632A3D6DABA1B069DE9459D15E58AE12130E2414DF92C36DCBDFE2EC3EB17E37393035ED810FBB857D971ECD41347B09C5C8DEEAB060E2759549A05C37A2C93F30CF906A9C59991DA921848363CEB06CF9914E76E1635AA0337A540470C9B3E58D152FE692AB3A1AB5F3E5C72598428DFB9D46E77C32001CC1E942902A4A1CD94D526042D3C16AE79A7F440F06ACC331E445E47FBCEA3AD5B2D4237E320C3DF1FD16CBA99AD93B136D971F4D7233898F1ED5E4017E4DE5B2243E6ADD776C4591E28B6F4A5FFA4AD7D273708D2C7C82BA28A0D621E9A10FAE863750C8FCBABCCF3F1D92E9E2FBD5D3D44B6C4C1A1A73C34523356A8B8DB1B8E7E6AF8B9A02FA03C705DEC578D6ECE7F1AB9C9498FFB1E283142B258342B53959B6E60BD23FDA24A53447049A6F5BD525B6E12DD60BEB5CC7BA0E245EDAEA2489AC0ACABCDBA4C6113F35ABFE30D69332BB6B05DD1430FE9A6AAC0AAE856F0391AC30814075085F8B784439EDD1BCF55FDFA0142424F7A9E0A92142AF3979C3D608D2CE99B9F63F9B3D487471F75D2C43FFBD137487DD9D9A8931D42992261E67FB1C531BC40500711FB83B2AA84C308AD061BE639698F3F2DFDB72864D950F0888A961261BCA7C0DBB78B9BDFB8024A51E3488D87AAEF8FD703A859E538886F0DE88A16AC90D2C596622E34E2E8D9685F918B6BE86AB5E3BD73194A21C9A4DB53FE0C88E027D8FB0621592BA8A8748267CE6EBEDFA75144E2DE1C1B39FB158095F9FEA12772216A718E4729E583B1516D8BDDF13736946073AA71E72F9AA068DD6C3E6D2C7D6BC66711B94BD75AD558DCDD77A1950096BB3922A482FD03B8ED9BA53DEC0083A8B2192848CEF5092D50FF687623A2ADDCBA7D5E9B15759DBB535B6C1ABA01CFB857BCADC6506F0F3E73DD649BC83A05FAA60CBED656F545732E30A838F95C7879D63077C18584E191E2F844D44FFD63C9223D61E38136856DFEF610BD812DA0B8E18FF2465A0FE9F4658AF94ED948B13B4E710AF03D3620";
    decaps_kats[0].msg = "8199CF923CE12126920108569C11CBF97CF03F44AF5CFA7D550E9B2AC7431982";
    decaps_kats[0].shared_key = "5D537CD0EF7B58F0FE95370473B96878F138ECC259ADFBF77EBD7328B822D9D9";

    // Iterate through KATs and validate
    foreach (decaps_kats[i]) begin
      parse_hex_to_array(decaps_kats[i].ek, kat_ek);
      parse_hex_to_array(decaps_kats[i].dk, kat_dk);
      parse_hex_to_array(decaps_kats[i].msg, kat_msg);
      parse_hex_to_array(decaps_kats[i].ciphertext, kat_ciphertext);
      parse_hex_to_array(decaps_kats[i].shared_key, kat_shared_key);

      `uvm_info("KAT", $sformatf("Running Decaps KAT %0d", i), UVM_LOW);

      // Wait for ready flag in MLKEM_STATUS
      ready = 0;
      while (!ready) begin
        reg_model.MLKEM_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", "Failed to read MLKEM_STATUS");
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("MLKEM_STATUS: %h", data), UVM_HIGH);
        end
        ready = data[0];
      end

      // Write MLKEM_DECAPS_KEY
      for(int j = 0; j < reg_model.MLKEM_DECAPS_KEY.m_mem.get_size(); j++) begin
        reg_model.MLKEM_DECAPS_KEY.m_mem.write(status, j, kat_dk[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLKEM_DECAPS_KEY[%0d]", i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLKEM_DECAPS_KEY[%0d]: %0h", j, kat_dk[j]), UVM_LOW);
        end
      end

      // Write MLKEM_CIPHERTEXT
      for(int j = 0; j < reg_model.MLKEM_CIPHERTEXT.m_mem.get_size(); j++) begin
        reg_model.MLKEM_CIPHERTEXT.m_mem.write(status, j, kat_ciphertext[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLKEM_CIPHERTEXT[%0d]", j));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLKEM_CIPHERTEXT[%0d]: %0h", j, kat_ciphertext[j]), UVM_LOW);
        end
      end

      // Trigger Decaps operation
      data = 'h00000003; // Decaps command
      reg_model.MLKEM_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE_FAIL", "Failed to write MLKEM_CTRL to trigger Decaps");
      end else begin
        `uvm_info("REG_WRITE_PASS", "Successfully wrote MLKEM_CTRL to trigger Decaps", UVM_LOW);
      end

      // Wait for ready flag in MLKEM_STATUS
      valid =0;
      while(!valid) begin
        reg_model.MLKEM_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end
      
      // Reading MLKEM_SHARED_KEY register
      foreach (reg_model.MLKEM_SHARED_KEY[j]) begin
        reg_model.MLKEM_SHARED_KEY[j].read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_SHARED_KEY[%0d]", j));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_SHARED_KEY[%0d]: %0h", j, data), UVM_LOW);
        end

        if (data !== kat_shared_key[j]) begin
          `uvm_error("VALIDATION_FAIL", $sformatf("SHARED KEY mismatch for KAT %0d at index %0d: Expected %h, Got %h", i, j, kat_shared_key[j], data));
        end else begin
          `uvm_info("VALIDATION_PASS", $sformatf("SHARED KEY match for KAT %0d at index %0d: %h", i, j, data), UVM_LOW);
        end
      end

      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end

    `uvm_info("KAT", $sformatf("Decaps KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



