// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
//======================================================================
//
// twiddle_rom.sv
// --------
// ROM contains twiddle factors for NTT and INTT
// 
//
//======================================================================

module ntt_twiddle_lookup 
    import ntt_defines_pkg::*;
#(
    parameter ADDR_WIDTH = 7,
    parameter DATA_WIDTH = 24
)
(

    input mode_t mode,
    input wire [ADDR_WIDTH-1:0] raddr,
    output logic [(3*DATA_WIDTH)-1:0] rdata
);

reg [(3*DATA_WIDTH)-1:0] ntt_twiddle_mem  [84:0];
reg [(3*DATA_WIDTH)-1:0] intt_twiddle_mem [84:0];

always_comb begin
    rdata = (mode == ct) ? ntt_twiddle_mem[raddr] : (mode inside {gs, pwm_intt}) ? intt_twiddle_mem[raddr] : 'h0;
end

logic [255 : 0][(DATA_WIDTH)-1:0] zeta;
logic [255 : 0][(DATA_WIDTH)-1:0] zetainv;

assign zeta[0] = 23'h000001;
assign zeta[1] = 23'h495E02;
assign zeta[2] = 23'h397567;
assign zeta[3] = 23'h396569;
assign zeta[4] = 23'h4F062B;
assign zeta[5] = 23'h53DF73;
assign zeta[6] = 23'h4FE033;
assign zeta[7] = 23'h4F066B;
assign zeta[8] = 23'h76B1AE;
assign zeta[9] = 23'h360DD5;
assign zeta[10] = 23'h28EDB0;
assign zeta[11] = 23'h207FE4;
assign zeta[12] = 23'h397283;
assign zeta[13] = 23'h70894A;
assign zeta[14] = 23'h088192;
assign zeta[15] = 23'h6D3DC8;
assign zeta[16] = 23'h4C7294;
assign zeta[17] = 23'h41E0B4;
assign zeta[18] = 23'h28A3D2;
assign zeta[19] = 23'h66528A;
assign zeta[20] = 23'h4A18A7;
assign zeta[21] = 23'h794034;
assign zeta[22] = 23'h0A52EE;
assign zeta[23] = 23'h6B7D81;
assign zeta[24] = 23'h4E9F1D;
assign zeta[25] = 23'h1A2877;
assign zeta[26] = 23'h2571DF;
assign zeta[27] = 23'h1649EE;
assign zeta[28] = 23'h7611BD;
assign zeta[29] = 23'h492BB7;
assign zeta[30] = 23'h2AF697;
assign zeta[31] = 23'h22D8D5;
assign zeta[32] = 23'h36F72A;
assign zeta[33] = 23'h30911E;
assign zeta[34] = 23'h29D13F;
assign zeta[35] = 23'h492673;
assign zeta[36] = 23'h50685F;
assign zeta[37] = 23'h2010A2;
assign zeta[38] = 23'h3887F7;
assign zeta[39] = 23'h11B2C3;
assign zeta[40] = 23'h0603A4;
assign zeta[41] = 23'h0E2BED;
assign zeta[42] = 23'h10B72C;
assign zeta[43] = 23'h4A5F35;
assign zeta[44] = 23'h1F9D15;
assign zeta[45] = 23'h428CD4;
assign zeta[46] = 23'h3177F4;
assign zeta[47] = 23'h20E612;
assign zeta[48] = 23'h341C1D;
assign zeta[49] = 23'h1AD873;
assign zeta[50] = 23'h736681;
assign zeta[51] = 23'h49553F;
assign zeta[52] = 23'h3952F6;
assign zeta[53] = 23'h62564A;
assign zeta[54] = 23'h65AD05;
assign zeta[55] = 23'h439A1C;
assign zeta[56] = 23'h53AA5F;
assign zeta[57] = 23'h30B622;
assign zeta[58] = 23'h087F38;
assign zeta[59] = 23'h3B0E6D;
assign zeta[60] = 23'h2C83DA;
assign zeta[61] = 23'h1C496E;
assign zeta[62] = 23'h330E2B;
assign zeta[63] = 23'h1C5B70;
assign zeta[64] = 23'h2EE3F1;
assign zeta[65] = 23'h137EB9;
assign zeta[66] = 23'h57A930;
assign zeta[67] = 23'h3AC6EF;
assign zeta[68] = 23'h3FD54C;
assign zeta[69] = 23'h4EB2EA;
assign zeta[70] = 23'h503EE1;
assign zeta[71] = 23'h7BB175;
assign zeta[72] = 23'h2648B4;
assign zeta[73] = 23'h1EF256;
assign zeta[74] = 23'h1D90A2;
assign zeta[75] = 23'h45A6D4;
assign zeta[76] = 23'h2AE59B;
assign zeta[77] = 23'h52589C;
assign zeta[78] = 23'h6EF1F5;
assign zeta[79] = 23'h3F7288;
assign zeta[80] = 23'h175102;
assign zeta[81] = 23'h075D59;
assign zeta[82] = 23'h1187BA;
assign zeta[83] = 23'h52ACA9;
assign zeta[84] = 23'h773E9E;
assign zeta[85] = 23'h0296D8;
assign zeta[86] = 23'h2592EC;
assign zeta[87] = 23'h4CFF12;
assign zeta[88] = 23'h404CE8;
assign zeta[89] = 23'h4AA582;
assign zeta[90] = 23'h1E54E6;
assign zeta[91] = 23'h4F16C1;
assign zeta[92] = 23'h1A7E79;
assign zeta[93] = 23'h03978F;
assign zeta[94] = 23'h4E4817;
assign zeta[95] = 23'h31B859;
assign zeta[96] = 23'h5884CC;
assign zeta[97] = 23'h1B4827;
assign zeta[98] = 23'h5B63D0;
assign zeta[99] = 23'h5D787A;
assign zeta[100] = 23'h35225E;
assign zeta[101] = 23'h400C7E;
assign zeta[102] = 23'h6C09D1;
assign zeta[103] = 23'h5BD532;
assign zeta[104] = 23'h6BC4D3;
assign zeta[105] = 23'h258ECB;
assign zeta[106] = 23'h2E534C;
assign zeta[107] = 23'h097A6C;
assign zeta[108] = 23'h3B8820;
assign zeta[109] = 23'h6D285C;
assign zeta[110] = 23'h2CA4F8;
assign zeta[111] = 23'h337CAA;
assign zeta[112] = 23'h14B2A0;
assign zeta[113] = 23'h558536;
assign zeta[114] = 23'h28F186;
assign zeta[115] = 23'h55795D;
assign zeta[116] = 23'h4AF670;
assign zeta[117] = 23'h234A86;
assign zeta[118] = 23'h75E826;
assign zeta[119] = 23'h78DE66;
assign zeta[120] = 23'h05528C;
assign zeta[121] = 23'h7ADF59;
assign zeta[122] = 23'h0F6E17;
assign zeta[123] = 23'h5BF3DA;
assign zeta[124] = 23'h459B7E;
assign zeta[125] = 23'h628B34;
assign zeta[126] = 23'h5DBECB;
assign zeta[127] = 23'h1A9E7B;
assign zeta[128] = 23'h0006D9;
assign zeta[129] = 23'h6257C5;
assign zeta[130] = 23'h574B3C;
assign zeta[131] = 23'h69A8EF;
assign zeta[132] = 23'h289838;
assign zeta[133] = 23'h64B5FE;
assign zeta[134] = 23'h7EF8F5;
assign zeta[135] = 23'h2A4E78;
assign zeta[136] = 23'h120A23;
assign zeta[137] = 23'h0154A8;
assign zeta[138] = 23'h09B7FF;
assign zeta[139] = 23'h435E87;
assign zeta[140] = 23'h437FF8;
assign zeta[141] = 23'h5CD5B4;
assign zeta[142] = 23'h4DC04E;
assign zeta[143] = 23'h4728AF;
assign zeta[144] = 23'h7F735D;
assign zeta[145] = 23'h0C8D0D;
assign zeta[146] = 23'h0F66D5;
assign zeta[147] = 23'h5A6D80;
assign zeta[148] = 23'h61AB98;
assign zeta[149] = 23'h185D96;
assign zeta[150] = 23'h437F31;
assign zeta[151] = 23'h468298;
assign zeta[152] = 23'h662960;
assign zeta[153] = 23'h4BD579;
assign zeta[154] = 23'h28DE06;
assign zeta[155] = 23'h465D8D;
assign zeta[156] = 23'h49B0E3;
assign zeta[157] = 23'h09B434;
assign zeta[158] = 23'h7C0DB3;
assign zeta[159] = 23'h5A68B0;
assign zeta[160] = 23'h409BA9;
assign zeta[161] = 23'h64D3D5;
assign zeta[162] = 23'h21762A;
assign zeta[163] = 23'h658591;
assign zeta[164] = 23'h246E39;
assign zeta[165] = 23'h48C39B;
assign zeta[166] = 23'h7BC759;
assign zeta[167] = 23'h4F5859;
assign zeta[168] = 23'h392DB2;
assign zeta[169] = 23'h230923;
assign zeta[170] = 23'h12EB67;
assign zeta[171] = 23'h454DF2;
assign zeta[172] = 23'h30C31C;
assign zeta[173] = 23'h285424;
assign zeta[174] = 23'h13232E;
assign zeta[175] = 23'h7FAF80;
assign zeta[176] = 23'h2DBFCB;
assign zeta[177] = 23'h022A0B;
assign zeta[178] = 23'h7E832C;
assign zeta[179] = 23'h26587A;
assign zeta[180] = 23'h6B3375;
assign zeta[181] = 23'h095B76;
assign zeta[182] = 23'h6BE1CC;
assign zeta[183] = 23'h5E061E;
assign zeta[184] = 23'h78E00D;
assign zeta[185] = 23'h628C37;
assign zeta[186] = 23'h3DA604;
assign zeta[187] = 23'h4AE53C;
assign zeta[188] = 23'h1F1D68;
assign zeta[189] = 23'h6330BB;
assign zeta[190] = 23'h7361B8;
assign zeta[191] = 23'h5EA06C;
assign zeta[192] = 23'h671AC7;
assign zeta[193] = 23'h201FC6;
assign zeta[194] = 23'h5BA4FF;
assign zeta[195] = 23'h60D772;
assign zeta[196] = 23'h08F201;
assign zeta[197] = 23'h6DE024;
assign zeta[198] = 23'h080E6D;
assign zeta[199] = 23'h56038E;
assign zeta[200] = 23'h695688;
assign zeta[201] = 23'h1E6D3E;
assign zeta[202] = 23'h2603BD;
assign zeta[203] = 23'h6A9DFA;
assign zeta[204] = 23'h07C017;
assign zeta[205] = 23'h6DBFD4;
assign zeta[206] = 23'h74D0BD;
assign zeta[207] = 23'h63E1E3;
assign zeta[208] = 23'h519573;
assign zeta[209] = 23'h7AB60D;
assign zeta[210] = 23'h2867BA;
assign zeta[211] = 23'h2DECD4;
assign zeta[212] = 23'h58018C;
assign zeta[213] = 23'h3F4CF5;
assign zeta[214] = 23'h0B7009;
assign zeta[215] = 23'h427E23;
assign zeta[216] = 23'h3CBD37;
assign zeta[217] = 23'h273333;
assign zeta[218] = 23'h673957;
assign zeta[219] = 23'h1A4B5D;
assign zeta[220] = 23'h196926;
assign zeta[221] = 23'h1EF206;
assign zeta[222] = 23'h11C14E;
assign zeta[223] = 23'h4C76C8;
assign zeta[224] = 23'h3CF42F;
assign zeta[225] = 23'h7FB19A;
assign zeta[226] = 23'h6AF66C;
assign zeta[227] = 23'h2E1669;
assign zeta[228] = 23'h3352D6;
assign zeta[229] = 23'h034760;
assign zeta[230] = 23'h085260;
assign zeta[231] = 23'h741E78;
assign zeta[232] = 23'h2F6316;
assign zeta[233] = 23'h6F0A11;
assign zeta[234] = 23'h07C0F1;
assign zeta[235] = 23'h776D0B;
assign zeta[236] = 23'h0D1FF0;
assign zeta[237] = 23'h345824;
assign zeta[238] = 23'h0223D4;
assign zeta[239] = 23'h68C559;
assign zeta[240] = 23'h5E8885;
assign zeta[241] = 23'h2FAA32;
assign zeta[242] = 23'h23FC65;
assign zeta[243] = 23'h5E6942;
assign zeta[244] = 23'h51E0ED;
assign zeta[245] = 23'h65ADB3;
assign zeta[246] = 23'h2CA5E6;
assign zeta[247] = 23'h79E1FE;
assign zeta[248] = 23'h7B4064;
assign zeta[249] = 23'h35E1DD;
assign zeta[250] = 23'h433AAC;
assign zeta[251] = 23'h464ADE;
assign zeta[252] = 23'h1CFE14;
assign zeta[253] = 23'h73F1CE;
assign zeta[254] = 23'h10170E;
assign zeta[255] = 23'h74B6D7;

//------------------------------------------------------------------------------------


assign zetainv[0] = 23'h7FE000;
assign zetainv[1] = 23'h3681FF;
assign zetainv[2] = 23'h466A9A;
assign zetainv[3] = 23'h467A98;
assign zetainv[4] = 23'h30D9D6;
assign zetainv[5] = 23'h2C008E;
assign zetainv[6] = 23'h2FFFCE;
assign zetainv[7] = 23'h30D996;
assign zetainv[8] = 23'h092E53;
assign zetainv[9] = 23'h49D22C;
assign zetainv[10] = 23'h56F251;
assign zetainv[11] = 23'h5F601D;
assign zetainv[12] = 23'h466D7E;
assign zetainv[13] = 23'h0F56B7;
assign zetainv[14] = 23'h775E6F;
assign zetainv[15] = 23'h12A239;
assign zetainv[16] = 23'h336D6D;
assign zetainv[17] = 23'h3DFF4D;
assign zetainv[18] = 23'h573C2F;
assign zetainv[19] = 23'h198D77;
assign zetainv[20] = 23'h35C75A;
assign zetainv[21] = 23'h069FCD;
assign zetainv[22] = 23'h758D13;
assign zetainv[23] = 23'h146280;
assign zetainv[24] = 23'h3140E4;
assign zetainv[25] = 23'h65B78A;
assign zetainv[26] = 23'h5A6E22;
assign zetainv[27] = 23'h699613;
assign zetainv[28] = 23'h09CE44;
assign zetainv[29] = 23'h36B44A;
assign zetainv[30] = 23'h54E96A;
assign zetainv[31] = 23'h5D072C;
assign zetainv[32] = 23'h48E8D7;
assign zetainv[33] = 23'h4F4EE3;
assign zetainv[34] = 23'h560EC2;
assign zetainv[35] = 23'h36B98E;
assign zetainv[36] = 23'h2F77A2;
assign zetainv[37] = 23'h5FCF5F;
assign zetainv[38] = 23'h47580A;
assign zetainv[39] = 23'h6E2D3E;
assign zetainv[40] = 23'h79DC5D;
assign zetainv[41] = 23'h71B414;
assign zetainv[42] = 23'h6F28D5;
assign zetainv[43] = 23'h3580CC;
assign zetainv[44] = 23'h6042EC;
assign zetainv[45] = 23'h3D532D;
assign zetainv[46] = 23'h4E680D;
assign zetainv[47] = 23'h5EF9EF;
assign zetainv[48] = 23'h4BC3E4;
assign zetainv[49] = 23'h65078E;
assign zetainv[50] = 23'h0C7980;
assign zetainv[51] = 23'h368AC2;
assign zetainv[52] = 23'h468D0B;
assign zetainv[53] = 23'h1D89B7;
assign zetainv[54] = 23'h1A32FC;
assign zetainv[55] = 23'h3C45E5;
assign zetainv[56] = 23'h2C35A2;
assign zetainv[57] = 23'h4F29DF;
assign zetainv[58] = 23'h7760C9;
assign zetainv[59] = 23'h44D194;
assign zetainv[60] = 23'h535C27;
assign zetainv[61] = 23'h639693;
assign zetainv[62] = 23'h4CD1D6;
assign zetainv[63] = 23'h638491;
assign zetainv[64] = 23'h50FC10;
assign zetainv[65] = 23'h6C6148;
assign zetainv[66] = 23'h2836D1;
assign zetainv[67] = 23'h451912;
assign zetainv[68] = 23'h400AB5;
assign zetainv[69] = 23'h312D17;
assign zetainv[70] = 23'h2FA120;
assign zetainv[71] = 23'h042E8C;
assign zetainv[72] = 23'h59974D;
assign zetainv[73] = 23'h60EDAB;
assign zetainv[74] = 23'h624F5F;
assign zetainv[75] = 23'h3A392D;
assign zetainv[76] = 23'h54FA66;
assign zetainv[77] = 23'h2D8765;
assign zetainv[78] = 23'h10EE0C;
assign zetainv[79] = 23'h406D79;
assign zetainv[80] = 23'h688EFF;
assign zetainv[81] = 23'h7882A8;
assign zetainv[82] = 23'h6E5847;
assign zetainv[83] = 23'h2D3358;
assign zetainv[84] = 23'h08A163;
assign zetainv[85] = 23'h7D4929;
assign zetainv[86] = 23'h5A4D15;
assign zetainv[87] = 23'h32E0EF;
assign zetainv[88] = 23'h3F9319;
assign zetainv[89] = 23'h353A7F;
assign zetainv[90] = 23'h618B1B;
assign zetainv[91] = 23'h30C940;
assign zetainv[92] = 23'h656188;
assign zetainv[93] = 23'h7C4872;
assign zetainv[94] = 23'h3197EA;
assign zetainv[95] = 23'h4E27A8;
assign zetainv[96] = 23'h275B35;
assign zetainv[97] = 23'h6497DA;
assign zetainv[98] = 23'h247C31;
assign zetainv[99] = 23'h226787;
assign zetainv[100] = 23'h4ABDA3;
assign zetainv[101] = 23'h3FD383;
assign zetainv[102] = 23'h13D630;
assign zetainv[103] = 23'h240ACF;
assign zetainv[104] = 23'h141B2E;
assign zetainv[105] = 23'h5A5136;
assign zetainv[106] = 23'h518CB5;
assign zetainv[107] = 23'h766595;
assign zetainv[108] = 23'h4457E1;
assign zetainv[109] = 23'h12B7A5;
assign zetainv[110] = 23'h533B09;
assign zetainv[111] = 23'h4C6357;
assign zetainv[112] = 23'h6B2D61;
assign zetainv[113] = 23'h2A5ACB;
assign zetainv[114] = 23'h56EE7B;
assign zetainv[115] = 23'h2A66A4;
assign zetainv[116] = 23'h34E991;
assign zetainv[117] = 23'h5C957B;
assign zetainv[118] = 23'h09F7DB;
assign zetainv[119] = 23'h07019B;
assign zetainv[120] = 23'h7A8D75;
assign zetainv[121] = 23'h0500A8;
assign zetainv[122] = 23'h7071EA;
assign zetainv[123] = 23'h23EC27;
assign zetainv[124] = 23'h3A4483;
assign zetainv[125] = 23'h1D54CD;
assign zetainv[126] = 23'h222136;
assign zetainv[127] = 23'h654186;
assign zetainv[128] = 23'h7FD928;
assign zetainv[129] = 23'h1D883C;
assign zetainv[130] = 23'h2894C5;
assign zetainv[131] = 23'h163712;
assign zetainv[132] = 23'h5747C9;
assign zetainv[133] = 23'h1B2A03;
assign zetainv[134] = 23'h00E70C;
assign zetainv[135] = 23'h559189;
assign zetainv[136] = 23'h6DD5DE;
assign zetainv[137] = 23'h7E8B59;
assign zetainv[138] = 23'h762802;
assign zetainv[139] = 23'h3C817A;
assign zetainv[140] = 23'h3C6009;
assign zetainv[141] = 23'h230A4D;
assign zetainv[142] = 23'h321FB3;
assign zetainv[143] = 23'h38B752;
assign zetainv[144] = 23'h006CA4;
assign zetainv[145] = 23'h7352F4;
assign zetainv[146] = 23'h70792C;
assign zetainv[147] = 23'h257281;
assign zetainv[148] = 23'h1E3469;
assign zetainv[149] = 23'h67826B;
assign zetainv[150] = 23'h3C60D0;
assign zetainv[151] = 23'h395D69;
assign zetainv[152] = 23'h19B6A1;
assign zetainv[153] = 23'h340A88;
assign zetainv[154] = 23'h5701FB;
assign zetainv[155] = 23'h398274;
assign zetainv[156] = 23'h362F1E;
assign zetainv[157] = 23'h762BCD;
assign zetainv[158] = 23'h03D24E;
assign zetainv[159] = 23'h257751;
assign zetainv[160] = 23'h3F4458;
assign zetainv[161] = 23'h1B0C2C;
assign zetainv[162] = 23'h5E69D7;
assign zetainv[163] = 23'h1A5A70;
assign zetainv[164] = 23'h5B71C8;
assign zetainv[165] = 23'h371C66;
assign zetainv[166] = 23'h0418A8;
assign zetainv[167] = 23'h3087A8;
assign zetainv[168] = 23'h46B24F;
assign zetainv[169] = 23'h5CD6DE;
assign zetainv[170] = 23'h6CF49A;
assign zetainv[171] = 23'h3A920F;
assign zetainv[172] = 23'h4F1CE5;
assign zetainv[173] = 23'h578BDD;
assign zetainv[174] = 23'h6CBCD3;
assign zetainv[175] = 23'h003081;
assign zetainv[176] = 23'h522036;
assign zetainv[177] = 23'h7DB5F6;
assign zetainv[178] = 23'h015CD5;
assign zetainv[179] = 23'h598787;
assign zetainv[180] = 23'h14AC8C;
assign zetainv[181] = 23'h76848B;
assign zetainv[182] = 23'h13FE35;
assign zetainv[183] = 23'h21D9E3;
assign zetainv[184] = 23'h06FFF4;
assign zetainv[185] = 23'h1D53CA;
assign zetainv[186] = 23'h4239FD;
assign zetainv[187] = 23'h34FAC5;
assign zetainv[188] = 23'h60C299;
assign zetainv[189] = 23'h1CAF46;
assign zetainv[190] = 23'h0C7E49;
assign zetainv[191] = 23'h213F95;
assign zetainv[192] = 23'h18C53A;
assign zetainv[193] = 23'h5FC03B;
assign zetainv[194] = 23'h243B02;
assign zetainv[195] = 23'h1F088F;
assign zetainv[196] = 23'h76EE00;
assign zetainv[197] = 23'h11FFDD;
assign zetainv[198] = 23'h77D194;
assign zetainv[199] = 23'h29DC73;
assign zetainv[200] = 23'h168979;
assign zetainv[201] = 23'h6172C3;
assign zetainv[202] = 23'h59DC44;
assign zetainv[203] = 23'h154207;
assign zetainv[204] = 23'h781FEA;
assign zetainv[205] = 23'h12202D;
assign zetainv[206] = 23'h0B0F44;
assign zetainv[207] = 23'h1BFE1E;
assign zetainv[208] = 23'h2E4A8E;
assign zetainv[209] = 23'h0529F4;
assign zetainv[210] = 23'h577847;
assign zetainv[211] = 23'h51F32D;
assign zetainv[212] = 23'h27DE75;
assign zetainv[213] = 23'h40930C;
assign zetainv[214] = 23'h746FF8;
assign zetainv[215] = 23'h3D61DE;
assign zetainv[216] = 23'h4322CA;
assign zetainv[217] = 23'h58ACCE;
assign zetainv[218] = 23'h18A6AA;
assign zetainv[219] = 23'h6594A4;
assign zetainv[220] = 23'h6676DB;
assign zetainv[221] = 23'h60EDFB;
assign zetainv[222] = 23'h6E1EB3;
assign zetainv[223] = 23'h336939;
assign zetainv[224] = 23'h42EBD2;
assign zetainv[225] = 23'h002E67;
assign zetainv[226] = 23'h14E995;
assign zetainv[227] = 23'h51C998;
assign zetainv[228] = 23'h4C8D2B;
assign zetainv[229] = 23'h7C98A1;
assign zetainv[230] = 23'h778DA1;
assign zetainv[231] = 23'h0BC189;
assign zetainv[232] = 23'h507CEB;
assign zetainv[233] = 23'h10D5F0;
assign zetainv[234] = 23'h781F10;
assign zetainv[235] = 23'h0872F6;
assign zetainv[236] = 23'h72C011;
assign zetainv[237] = 23'h4B87DD;
assign zetainv[238] = 23'h7DBC2D;
assign zetainv[239] = 23'h171AA8;
assign zetainv[240] = 23'h21577C;
assign zetainv[241] = 23'h5035CF;
assign zetainv[242] = 23'h5BE39C;
assign zetainv[243] = 23'h2176BF;
assign zetainv[244] = 23'h2DFF14;
assign zetainv[245] = 23'h1A324E;
assign zetainv[246] = 23'h533A1B;
assign zetainv[247] = 23'h05FE03;
assign zetainv[248] = 23'h049F9D;
assign zetainv[249] = 23'h49FE24;
assign zetainv[250] = 23'h3CA555;
assign zetainv[251] = 23'h399523;
assign zetainv[252] = 23'h62E1ED;
assign zetainv[253] = 23'h0BEE33;
assign zetainv[254] = 23'h6FC8F3;
assign zetainv[255] = 23'h0B292A;

// assign ntt_twiddle_mem[0]  = 'h000001;
assign ntt_twiddle_mem[0]  = {zeta[3],  zeta[2],  zeta[1]};
assign ntt_twiddle_mem[1]  = {zeta[9],  zeta[8],  zeta[4]};
assign ntt_twiddle_mem[2]  = {zeta[11], zeta[10], zeta[5]};
assign ntt_twiddle_mem[3]  = {zeta[13], zeta[12], zeta[6]};
assign ntt_twiddle_mem[4]  = {zeta[15], zeta[14], zeta[7]};
assign ntt_twiddle_mem[5]  = {zeta[33], zeta[32], zeta[16]};
assign ntt_twiddle_mem[6]  = {zeta[35], zeta[34], zeta[17]};
assign ntt_twiddle_mem[7]  = {zeta[37], zeta[36], zeta[18]};
assign ntt_twiddle_mem[8]  = {zeta[39], zeta[38], zeta[19]};
assign ntt_twiddle_mem[9]  = {zeta[41], zeta[40], zeta[20]};
assign ntt_twiddle_mem[10] = {zeta[43], zeta[42], zeta[21]};
assign ntt_twiddle_mem[11] = {zeta[45], zeta[44], zeta[22]};
assign ntt_twiddle_mem[12] = {zeta[47], zeta[46], zeta[23]};
assign ntt_twiddle_mem[13] = {zeta[49], zeta[48], zeta[24]};
assign ntt_twiddle_mem[14] = {zeta[51], zeta[50], zeta[25]};
assign ntt_twiddle_mem[15] = {zeta[53], zeta[52], zeta[26]};
assign ntt_twiddle_mem[16] = {zeta[55], zeta[54], zeta[27]};
assign ntt_twiddle_mem[17] = {zeta[57], zeta[56], zeta[28]};
assign ntt_twiddle_mem[18] = {zeta[59], zeta[58], zeta[29]};
assign ntt_twiddle_mem[19] = {zeta[61], zeta[60], zeta[30]};
assign ntt_twiddle_mem[20] = {zeta[63], zeta[62], zeta[31]};
assign ntt_twiddle_mem[21] = {zeta[129], zeta[128], zeta[64]};
assign ntt_twiddle_mem[22] = {zeta[131], zeta[130], zeta[65]};
assign ntt_twiddle_mem[23] = {zeta[133], zeta[132], zeta[66]};
assign ntt_twiddle_mem[24] = {zeta[135], zeta[134], zeta[67]};
assign ntt_twiddle_mem[25] = {zeta[137], zeta[136], zeta[68]};
assign ntt_twiddle_mem[26] = {zeta[139], zeta[138], zeta[69]};
assign ntt_twiddle_mem[27] = {zeta[141], zeta[140], zeta[70]};
assign ntt_twiddle_mem[28] = {zeta[143], zeta[142], zeta[71]};
assign ntt_twiddle_mem[29] = {zeta[145], zeta[144], zeta[72]};
assign ntt_twiddle_mem[30] = {zeta[147], zeta[146], zeta[73]};
assign ntt_twiddle_mem[31] = {zeta[149], zeta[148], zeta[74]};
assign ntt_twiddle_mem[32] = {zeta[151], zeta[150], zeta[75]};
assign ntt_twiddle_mem[33] = {zeta[153], zeta[152], zeta[76]};
assign ntt_twiddle_mem[34] = {zeta[155], zeta[154], zeta[77]};
assign ntt_twiddle_mem[35] = {zeta[157], zeta[156], zeta[78]};
assign ntt_twiddle_mem[36] = {zeta[159], zeta[158], zeta[79]};
assign ntt_twiddle_mem[37] = {zeta[161], zeta[160], zeta[80]};
assign ntt_twiddle_mem[38] = {zeta[163], zeta[162], zeta[81]};
assign ntt_twiddle_mem[39] = {zeta[165], zeta[164], zeta[82]};
assign ntt_twiddle_mem[40] = {zeta[167], zeta[166], zeta[83]};
assign ntt_twiddle_mem[41] = {zeta[169], zeta[168], zeta[84]};
assign ntt_twiddle_mem[42] = {zeta[171], zeta[170], zeta[85]};
assign ntt_twiddle_mem[43] = {zeta[173], zeta[172], zeta[86]};
assign ntt_twiddle_mem[44] = {zeta[175], zeta[174], zeta[87]};
assign ntt_twiddle_mem[45] = {zeta[177], zeta[176], zeta[88]};
assign ntt_twiddle_mem[46] = {zeta[179], zeta[178], zeta[89]};
assign ntt_twiddle_mem[47] = {zeta[181], zeta[180], zeta[90]};
assign ntt_twiddle_mem[48] = {zeta[183], zeta[182], zeta[91]};
assign ntt_twiddle_mem[49] = {zeta[185], zeta[184], zeta[92]};
assign ntt_twiddle_mem[50] = {zeta[187], zeta[186], zeta[93]};
assign ntt_twiddle_mem[51] = {zeta[189], zeta[188], zeta[94]};
assign ntt_twiddle_mem[52] = {zeta[191], zeta[190], zeta[95]};
assign ntt_twiddle_mem[53] = {zeta[193], zeta[192], zeta[96]};
assign ntt_twiddle_mem[54] = {zeta[195], zeta[194], zeta[97]};
assign ntt_twiddle_mem[55] = {zeta[197], zeta[196], zeta[98]};
assign ntt_twiddle_mem[56] = {zeta[199], zeta[198], zeta[99]};
assign ntt_twiddle_mem[57] = {zeta[201], zeta[200], zeta[100]};
assign ntt_twiddle_mem[58] = {zeta[203], zeta[202], zeta[101]};
assign ntt_twiddle_mem[59] = {zeta[205], zeta[204], zeta[102]};
assign ntt_twiddle_mem[60] = {zeta[207], zeta[206], zeta[103]};
assign ntt_twiddle_mem[61] = {zeta[209], zeta[208], zeta[104]};
assign ntt_twiddle_mem[62] = {zeta[211], zeta[210], zeta[105]};
assign ntt_twiddle_mem[63] = {zeta[213], zeta[212], zeta[106]};
assign ntt_twiddle_mem[64] = {zeta[215], zeta[214], zeta[107]};
assign ntt_twiddle_mem[65] = {zeta[217], zeta[216], zeta[108]};
assign ntt_twiddle_mem[66] = {zeta[219], zeta[218], zeta[109]};
assign ntt_twiddle_mem[67] = {zeta[221], zeta[220], zeta[110]};
assign ntt_twiddle_mem[68] = {zeta[223], zeta[222], zeta[111]};
assign ntt_twiddle_mem[69] = {zeta[225], zeta[224], zeta[112]};
assign ntt_twiddle_mem[70] = {zeta[227], zeta[226], zeta[113]};
assign ntt_twiddle_mem[71] = {zeta[229], zeta[228], zeta[114]};
assign ntt_twiddle_mem[72] = {zeta[231], zeta[230], zeta[115]};
assign ntt_twiddle_mem[73] = {zeta[233], zeta[232], zeta[116]};
assign ntt_twiddle_mem[74] = {zeta[235], zeta[234], zeta[117]};
assign ntt_twiddle_mem[75] = {zeta[237], zeta[236], zeta[118]};
assign ntt_twiddle_mem[76] = {zeta[239], zeta[238], zeta[119]};
assign ntt_twiddle_mem[77] = {zeta[241], zeta[240], zeta[120]};
assign ntt_twiddle_mem[78] = {zeta[243], zeta[242], zeta[121]};
assign ntt_twiddle_mem[79] = {zeta[245], zeta[244], zeta[122]};
assign ntt_twiddle_mem[80] = {zeta[247], zeta[246], zeta[123]};
assign ntt_twiddle_mem[81] = {zeta[249], zeta[248], zeta[124]};
assign ntt_twiddle_mem[82] = {zeta[251], zeta[250], zeta[125]};
assign ntt_twiddle_mem[83] = {zeta[253], zeta[252], zeta[126]};
assign ntt_twiddle_mem[84] = {zeta[255], zeta[254], zeta[127]};
//--------------------------------------------------------

assign intt_twiddle_mem[0]  = {zetainv[127], zetainv[254], zetainv[255]};
assign intt_twiddle_mem[1]  = {zetainv[126], zetainv[252], zetainv[253]};
assign intt_twiddle_mem[2]  = {zetainv[125], zetainv[250], zetainv[251]};
assign intt_twiddle_mem[3]  = {zetainv[124], zetainv[248], zetainv[249]};
assign intt_twiddle_mem[4]  = {zetainv[123], zetainv[246], zetainv[247]};
assign intt_twiddle_mem[5]  = {zetainv[122], zetainv[244], zetainv[245]};
assign intt_twiddle_mem[6]  = {zetainv[121], zetainv[242], zetainv[243]};
assign intt_twiddle_mem[7]  = {zetainv[120], zetainv[240], zetainv[241]};
assign intt_twiddle_mem[8]  = {zetainv[119], zetainv[238], zetainv[239]};
assign intt_twiddle_mem[9]  = {zetainv[118], zetainv[236], zetainv[237]};
assign intt_twiddle_mem[10] = {zetainv[117], zetainv[234], zetainv[235]};
assign intt_twiddle_mem[11] = {zetainv[116], zetainv[232], zetainv[233]};
assign intt_twiddle_mem[12] = {zetainv[115], zetainv[230], zetainv[231]};
assign intt_twiddle_mem[13] = {zetainv[114], zetainv[228], zetainv[229]};
assign intt_twiddle_mem[14] = {zetainv[113], zetainv[226], zetainv[227]};
assign intt_twiddle_mem[15] = {zetainv[112], zetainv[224], zetainv[225]};
assign intt_twiddle_mem[16] = {zetainv[111], zetainv[222], zetainv[223]};
assign intt_twiddle_mem[17] = {zetainv[110], zetainv[220], zetainv[221]};
assign intt_twiddle_mem[18] = {zetainv[109], zetainv[218], zetainv[219]};
assign intt_twiddle_mem[19] = {zetainv[108], zetainv[216], zetainv[217]};
assign intt_twiddle_mem[20] = {zetainv[107], zetainv[214], zetainv[215]};
assign intt_twiddle_mem[21] = {zetainv[106], zetainv[212], zetainv[213]};
assign intt_twiddle_mem[22] = {zetainv[105], zetainv[210], zetainv[211]};
assign intt_twiddle_mem[23] = {zetainv[104], zetainv[208], zetainv[209]};
assign intt_twiddle_mem[24] = {zetainv[103], zetainv[206], zetainv[207]};
assign intt_twiddle_mem[25] = {zetainv[102], zetainv[204], zetainv[205]};
assign intt_twiddle_mem[26] = {zetainv[101], zetainv[202], zetainv[203]};
assign intt_twiddle_mem[27] = {zetainv[100], zetainv[200], zetainv[201]};
assign intt_twiddle_mem[28] = {zetainv[99], zetainv[198], zetainv[199]};
assign intt_twiddle_mem[29] = {zetainv[98], zetainv[196], zetainv[197]};
assign intt_twiddle_mem[30] = {zetainv[97], zetainv[194], zetainv[195]};
assign intt_twiddle_mem[31] = {zetainv[96], zetainv[192], zetainv[193]};
assign intt_twiddle_mem[32] = {zetainv[95], zetainv[190], zetainv[191]};
assign intt_twiddle_mem[33] = {zetainv[94], zetainv[188], zetainv[189]};
assign intt_twiddle_mem[34] = {zetainv[93], zetainv[186], zetainv[187]};
assign intt_twiddle_mem[35] = {zetainv[92], zetainv[184], zetainv[185]};
assign intt_twiddle_mem[36] = {zetainv[91], zetainv[182], zetainv[183]};
assign intt_twiddle_mem[37] = {zetainv[90], zetainv[180], zetainv[181]};
assign intt_twiddle_mem[38] = {zetainv[89], zetainv[178], zetainv[179]};
assign intt_twiddle_mem[39] = {zetainv[88], zetainv[176], zetainv[177]};
assign intt_twiddle_mem[40] = {zetainv[87], zetainv[174], zetainv[175]};
assign intt_twiddle_mem[41] = {zetainv[86], zetainv[172], zetainv[173]};
assign intt_twiddle_mem[42] = {zetainv[85], zetainv[170], zetainv[171]};
assign intt_twiddle_mem[43] = {zetainv[84], zetainv[168], zetainv[169]};
assign intt_twiddle_mem[44] = {zetainv[83], zetainv[166], zetainv[167]};
assign intt_twiddle_mem[45] = {zetainv[82], zetainv[164], zetainv[165]};
assign intt_twiddle_mem[46] = {zetainv[81], zetainv[162], zetainv[163]};
assign intt_twiddle_mem[47] = {zetainv[80], zetainv[160], zetainv[161]};
assign intt_twiddle_mem[48] = {zetainv[79], zetainv[158], zetainv[159]};
assign intt_twiddle_mem[49] = {zetainv[78], zetainv[156], zetainv[157]};
assign intt_twiddle_mem[50] = {zetainv[77], zetainv[154], zetainv[155]};
assign intt_twiddle_mem[51] = {zetainv[76], zetainv[152], zetainv[153]};
assign intt_twiddle_mem[52] = {zetainv[75], zetainv[150], zetainv[151]};
assign intt_twiddle_mem[53] = {zetainv[74], zetainv[148], zetainv[149]};
assign intt_twiddle_mem[54] = {zetainv[73], zetainv[146], zetainv[147]};
assign intt_twiddle_mem[55] = {zetainv[72], zetainv[144], zetainv[145]};
assign intt_twiddle_mem[56] = {zetainv[71], zetainv[142], zetainv[143]};
assign intt_twiddle_mem[57] = {zetainv[70], zetainv[140], zetainv[141]};
assign intt_twiddle_mem[58] = {zetainv[69], zetainv[138], zetainv[139]};
assign intt_twiddle_mem[59] = {zetainv[68], zetainv[136], zetainv[137]};
assign intt_twiddle_mem[60] = {zetainv[67], zetainv[134], zetainv[135]};
assign intt_twiddle_mem[61] = {zetainv[66], zetainv[132], zetainv[133]};
assign intt_twiddle_mem[62] = {zetainv[65], zetainv[130], zetainv[131]};
assign intt_twiddle_mem[63] = {zetainv[64], zetainv[128], zetainv[129]};
assign intt_twiddle_mem[64] = {zetainv[31], zetainv[62], zetainv[63]};
assign intt_twiddle_mem[65] = {zetainv[30], zetainv[60], zetainv[61]};
assign intt_twiddle_mem[66] = {zetainv[29], zetainv[58], zetainv[59]}; 
assign intt_twiddle_mem[67] = {zetainv[28], zetainv[56], zetainv[57]};
assign intt_twiddle_mem[68] = {zetainv[27], zetainv[54], zetainv[55]};
assign intt_twiddle_mem[69] = {zetainv[26], zetainv[52], zetainv[53]};
assign intt_twiddle_mem[70] = {zetainv[25], zetainv[50], zetainv[51]};
assign intt_twiddle_mem[71] = {zetainv[24], zetainv[48], zetainv[49]};
assign intt_twiddle_mem[72] = {zetainv[23], zetainv[46], zetainv[47]};
assign intt_twiddle_mem[73] = {zetainv[22], zetainv[44], zetainv[45]};
assign intt_twiddle_mem[74] = {zetainv[21], zetainv[42], zetainv[43]};
assign intt_twiddle_mem[75] = {zetainv[20], zetainv[40], zetainv[41]};
assign intt_twiddle_mem[76] = {zetainv[19], zetainv[38], zetainv[39]};
assign intt_twiddle_mem[77] = {zetainv[18], zetainv[36], zetainv[37]};
assign intt_twiddle_mem[78] = {zetainv[17], zetainv[34], zetainv[35]};
assign intt_twiddle_mem[79] = {zetainv[16], zetainv[32], zetainv[33]};
assign intt_twiddle_mem[80] = {zetainv[7], zetainv[14], zetainv[15]};
assign intt_twiddle_mem[81] = {zetainv[6], zetainv[12], zetainv[13]};
assign intt_twiddle_mem[82] = {zetainv[5], zetainv[10], zetainv[11]};
assign intt_twiddle_mem[83] = {zetainv[4], zetainv[8], zetainv[9]};
assign intt_twiddle_mem[84] = {zetainv[1], zetainv[2], zetainv[3]};


endmodule