//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef struct {
  string seed_d;       // Input SEED_D
  string seed_z;       // Input SEED_Z
  string expected_PK;  // Expected Public Key
  string expected_SK;  // Expected Secret Key
} mlkem_keygen_kat_t;

class ML_KEM_keygen_KATs_sequence extends mldsa_bench_sequence_base;

  `uvm_object_utils(ML_KEM_keygen_KATs_sequence);

    
    // KAT arrays
  mlkem_keygen_kat_t keygen_kats[];
  bit [31:0] kat_seed_d [];
  bit [31:0] kat_seed_z [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    keygen_kats = new[1];
    kat_seed_d = new[8];
    kat_seed_z = new[8];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // KeyGen KATs
    keygen_kats[0].seed_z = "0A064D6C06CEAB73E59CFCA9FF6402255A326AEF1E9CB678BF36929DAFE29A58";
    keygen_kats[0].seed_d = "2B5330C4F23BFDFD5C31F050BA3B38235324BF032372FC12D04DD08920F0BD59";
    keygen_kats[0].expected_PK = "B24174A5B00DBF520CB9E3783D482E03CA3166D40D082A7BAB664845B617ADD98C07C6A3C3204F812035683A1D4F10AC1DE764706CCE96D75832A462A8B1B82CF471CBF808A26508D9FAA543F2CD980377D6F794367938064B6DD388C529756963B12CA594B306AB3F0EBBB6ED47601AEC1074A2B0D1B41717F8C695F174EF734052077E53DC9F47316B6608B7EDB54EA3631A36BB8D842CAF27367C15C18DDBA7AFE62AA572133384CB872555948A165F204C2CB4503C9D8ACE5F5217194A67EBD2A72F99562F98B2B773B6965C071BF11DEED395BC153ED6967492D88D5EF32D05E008B7958A2F36B9DB06CCDC52A626417966B19C5079A9892BA426A0362FB18E7EC07FFDC0C5DBE264DEEC41BC83A573599A25A8909B2476682336CEC9A396201A000A9C1BE792D9988FBC03C24855C1B242AE27A127CD36415CFB0D98CCBB9BD83AF5988D743773ACEA4201AC935E7CCC46E92D8E84A9D70CC626965429450980E0782EE11CD91169CE94BF89C14EC10B900EB4B77129A859039AD1253E5657B261E9855BC4B0F504C478D58F4A388215A0715168109526C2DAC555007C66E10B79EB92471ACC9A640805BD947EEA45B66A2C02D5B7C9029945B581666D470CD2654EB51C3304AC52CB11382B8628553B63742C41B293467B754DF8F52A7B9A5EF2359BF34025A9318DF92B1471EC529E895814999C551356ECC9CA945641067B16AC04B4169CC2F8A3B9A005047AC1AA4DF27FF284C7AB19A800629B5A85B06834623AC018D2E4CA1CA197D7B458C185BE0BA9B4703811F8628D13B690602544BD69AFAE215F5BDB51315CB570D48D8B55120D50560E59594C8B5603FBCC7E484EAF591070865FADD495C4D67BFC67CF1CB94ACD50C8970A226C0BC0FFA186BDC51DD235AC8D085F348374C88C6206E147233104306916E30635F0AB1B956644E02A4EE2BCC3246088D3D570A617A63150B32BD50DAA555DD6BB8B6D34C0CBA83A41C23B48B39708D7578D33C5A60AA28430CB10BA264D158ABFF301A00732BD95539190436AD02F89315CE921499C04305D81CFB7997ABA4B2D65639A34901B67972C9A2355B5A10E91F955E0A95FF33A21FA4A8B8E018EA6E43F34462DAF95A29DCC719C2B7EEAE50350497006F6AC53D28FCBF90845B02A8846C58D6494C0C603283476AF121767A9600C83A9E92B8D7B19C2680B1948044B807C9EA7EC94BE30CF3AEA676D16159FA3BC97C055ED0A439AF5C2F085BC0680A5DED6820843C3D3F65138E5ACE48C7A0C11037161674826084FD9BA3113223F18564A9B8DD98472D1837AB85B66E2C2638A4A8D9DD6C361BA6B86629FED9B6E76DC75B258908B750117E8A4763A1C0C0BBE5E2616C5D55B60720371F06D63893061FA6B3C76A600179B52F0C319F47A10189A0F566A7292C40CD9980C0112F265660C3B4F60736A9693454A7B861F834D35B838F8A647771630BCBC1F23F6AA887CB6CBD582CC2240CDBA864167506A43C434C27EAD754484D232A83BC40C2218306816030A20765A5470217E5B2C90846344CD8BC2C498B770E83CD1959DC152BCCB4ACEAB36ABF7F3618C1247F5DB201310C0A1E574FA547C398CC5A44AC23685B64D07B8F6614016C4271B71C650A8B520A5AFA08BA04EE51646B8A7FB652D3AF57A4010558F856FACC9911E09B332C5870EDB61E8E850BB1949AE5755C1FBA2CC472073029FD6542BCDA71B7952BCF811608F2A88291A04F2664BB1112E27B1235B16C19203214E79145A318C5110152DA36BB21ACA73801185D6B8B1F6A344B33B3E550FB5DC29BCD19846E84074BBC8F7580CD347B52F12A7D1616C55A2CD1F5C4AA86702DD530FA05A641302A16127468E85522E567570B65FC3F834D85A20973A0EB2B210D5812CFDFB881CC3AA06AB4CB77BBA7CDC6BCEE53C020B3343B9BD9A8298AD2055EE1A6070849140A86288721815C79734773F4097CF4741CC9635A30C8100B20733D3980B350393FAAC4CD0E66E4737C681DBBCC8D7953FA77454C422AD870E278B1121C33C8273370E5B686A6AAB17FCA3B67A3040D6491241BF5E3072FBDC1E422413FA5B4E9EE91EB3C936E21A5C7856942F44A55670A688A69E91A9A80BF4094C301DF705334DACB0CD929473829F34F37947D22B55C062F4CCF703EE3C1CC0BA7316DD658E6B6E0815F8FC9A70B1BBA325EC32E2930916";
    keygen_kats[0].expected_SK = "F7517C1258A61E1936F15B11DBBB33A7F7733CCCB2D9493CBF29945C751E2519347AA3894541CC2F1010D590447872547238C2FDEA5764BA0D098030962A0EC6BB816B077FF4EC2EF1E6B4AB45B21DC99EA433B4B8F4CB36A41D1497A06BDC43CB79AA0F739E6286AFA063B908138FE837330E48A47A097EFADC3AACBAA059B320B2B81DAD5A9C27B24A66D74B3AAB48E6E355AAF18074DA3E9BE2418CC143388153DF649572036ABCA2096C85839E034D34FCA6B9530B07E80534479A3BB6B7B09922FB4058A20B2585A74C45C14FFE076BF8D40CF5C922E14A3D34325B5909729C870B36BCC17964590E51CCDE66B1425ACFAFBC5CECD10FB168005C04C65654B7574150F18C2362F18136A09CF12029BA371E008029B4B631021A252E756E3BC40E41030A3A2A52205A917EF4B0A66A8279A8B67309A2D35460085BBE18F221BB72409F004A894BA1AE2A31141389FB963DB3F0C0DA0A179FA30926DA2D817AA6FFF02BF656716AA87F7273B747741CBAB3ACFC112D3942C193DC32A31A2A0425854206B51807C960D93D6E361A5F29A6F15A417FD01D25E264C322C8696369FF5397EDC52D6D388BBAD6206729BA14D7855DF4424AE9C48AD11A19AAA2F8FBBE50BB6AC1208385E80C740C916AB540504758F7879B0D0B5B36C0053E564E15017E563966EF0162966B0A6A330A4079C9D01A89B43893E38C4064A247B1F98627EAAB80A1603A43C01FFC5D63DCA4DAEA501379CAAFF77BBF0C238B091318548168F4033B83A2D2C6026AD2973BA43C01914B27DC248805C762D980E7B427252B222DE59698BAAD02936E1135704CF80F531C13FB9828D1199762794B69762BFA3134BCA20AD4F799CE0B5F27586654D981598172E191B4B556457B27C1CDE17B2A9A4752466439693622C68DF2608CA84B86BC553CCCAB9D9C842387B8764C946917E26409DA1C92122273AB6124784D8B1475287A3492E2A90D770BDD116BF0FC0460C56A07D86DB686983A052D7E01392C5B34F8DB41D339808D2A9AEF44C845A6B67688AB74FB1218E7AF9D172DE406BE0A32CB40710FC33098B82A21AA719124EA3D12A28E87043AFE9B56CDC58534BB38E497512CB939CC3CB4D7D3ADFB2C9F4DB11100D76A77BB2CFAD308F3171AD0478411009B11E964D1721A1225A90A285073445B9E389F72B46AACF08EC5DB33F7E038D4CB4C8FF023A5D8BBFD543BED672ED38927807B285B0C3635A1BF554729EA595595C1A1718122821C446E72BA7C5C95F3CAB365B27CE4A283C745386F260320F56815A9704F4C2718D89F60754BD65434A65063665B723033AD8E2213B1562EC9296A370B0C8D5497691718BFFA1F65E26B3709B7A632945B592FBEA90588B0BEF3877630212DFE76792B40A0B4E173161AA641119FAF78905A7C3E59E3686A0B1654E48AB9C22D18BCA456D553DAB3436EE677AB7AB9ECE7416B7A90921A8742A9269742616BF22572A2C8FABBAFCCD1441E87C9AB64593AE50A5C9564834A08851462AFA41A3DB586D49835CBB8A5CF5950B85ABE5D1A64F8C82129AC488000474E5386B3429ADE528345582A8185010DC39D0DA6873D29BEBF3954A56902AC623ED9577103164A839B89BE158CA639C1EF483902A3A1AB1513CCEB62DEF158D0078593321EFFA057B0A17C854956A73C48D55C3B1511C4B43316C95C18FB784452DC4D2C904D30206F17B4644A755344462A034C3D55F04DE42843CAD248E256C2616A98D61024B1D9547C86B37625484C3373E0B786B1220C7EC1A3E75715277C014AC81FFC7A80135B90A9D65DFBDCB03050756ADC26949B1644BBA4EFF133BECB67FBA996C4958DC49C5824B8824433AECBE468DBFB3D46289F65B6528204BE31A8A22B828EA30766CE086E380A6A94EC119C3AC9005D2B8BE47AF0FA2E7C008B06C7CA9827B7E6A247A75717954726E4D96EC82B7EBD469F9C646612C2A785EC3EF1CB5CD5A76F7D006418B19FB3C8254A381320984D03F62244C72A55AA19F60A63EE0B900BA56287235D1D480E752AC905A57D3C99B7C3210E103C50FEC53E430926CC108F0240CE4E3A5116645B5BE79F03AC0D378B00FDA6206C5C5CBC551851243E8EAC7C7B28AA13592FF38065D6F8B73A66812AA415CE44162476008288AFAF1A02B24174A5B00DBF520CB9E3783D482E03CA3166D40D082A7BAB664845B617ADD98C07C6A3C3204F812035683A1D4F10AC1DE764706CCE96D75832A462A8B1B82CF471CBF808A26508D9FAA543F2CD980377D6F794367938064B6DD388C529756963B12CA594B306AB3F0EBBB6ED47601AEC1074A2B0D1B41717F8C695F174EF734052077E53DC9F47316B6608B7EDB54EA3631A36BB8D842CAF27367C15C18DDBA7AFE62AA572133384CB872555948A165F204C2CB4503C9D8ACE5F5217194A67EBD2A72F99562F98B2B773B6965C071BF11DEED395BC153ED6967492D88D5EF32D05E008B7958A2F36B9DB06CCDC52A626417966B19C5079A9892BA426A0362FB18E7EC07FFDC0C5DBE264DEEC41BC83A573599A25A8909B2476682336CEC9A396201A000A9C1BE792D9988FBC03C24855C1B242AE27A127CD36415CFB0D98CCBB9BD83AF5988D743773ACEA4201AC935E7CCC46E92D8E84A9D70CC626965429450980E0782EE11CD91169CE94BF89C14EC10B900EB4B77129A859039AD1253E5657B261E9855BC4B0F504C478D58F4A388215A0715168109526C2DAC555007C66E10B79EB92471ACC9A640805BD947EEA45B66A2C02D5B7C9029945B581666D470CD2654EB51C3304AC52CB11382B8628553B63742C41B293467B754DF8F52A7B9A5EF2359BF34025A9318DF92B1471EC529E895814999C551356ECC9CA945641067B16AC04B4169CC2F8A3B9A005047AC1AA4DF27FF284C7AB19A800629B5A85B06834623AC018D2E4CA1CA197D7B458C185BE0BA9B4703811F8628D13B690602544BD69AFAE215F5BDB51315CB570D48D8B55120D50560E59594C8B5603FBCC7E484EAF591070865FADD495C4D67BFC67CF1CB94ACD50C8970A226C0BC0FFA186BDC51DD235AC8D085F348374C88C6206E147233104306916E30635F0AB1B956644E02A4EE2BCC3246088D3D570A617A63150B32BD50DAA555DD6BB8B6D34C0CBA83A41C23B48B39708D7578D33C5A60AA28430CB10BA264D158ABFF301A00732BD95539190436AD02F89315CE921499C04305D81CFB7997ABA4B2D65639A34901B67972C9A2355B5A10E91F955E0A95FF33A21FA4A8B8E018EA6E43F34462DAF95A29DCC719C2B7EEAE50350497006F6AC53D28FCBF90845B02A8846C58D6494C0C603283476AF121767A9600C83A9E92B8D7B19C2680B1948044B807C9EA7EC94BE30CF3AEA676D16159FA3BC97C055ED0A439AF5C2F085BC0680A5DED6820843C3D3F65138E5ACE48C7A0C11037161674826084FD9BA3113223F18564A9B8DD98472D1837AB85B66E2C2638A4A8D9DD6C361BA6B86629FED9B6E76DC75B258908B750117E8A4763A1C0C0BBE5E2616C5D55B60720371F06D63893061FA6B3C76A600179B52F0C319F47A10189A0F566A7292C40CD9980C0112F265660C3B4F60736A9693454A7B861F834D35B838F8A647771630BCBC1F23F6AA887CB6CBD582CC2240CDBA864167506A43C434C27EAD754484D232A83BC40C2218306816030A20765A5470217E5B2C90846344CD8BC2C498B770E83CD1959DC152BCCB4ACEAB36ABF7F3618C1247F5DB201310C0A1E574FA547C398CC5A44AC23685B64D07B8F6614016C4271B71C650A8B520A5AFA08BA04EE51646B8A7FB652D3AF57A4010558F856FACC9911E09B332C5870EDB61E8E850BB1949AE5755C1FBA2CC472073029FD6542BCDA71B7952BCF811608F2A88291A04F2664BB1112E27B1235B16C19203214E79145A318C5110152DA36BB21ACA73801185D6B8B1F6A344B33B3E550FB5DC29BCD19846E84074BBC8F7580CD347B52F12A7D1616C55A2CD1F5C4AA86702DD530FA05A641302A16127468E85522E567570B65FC3F834D85A20973A0EB2B210D5812CFDFB881CC3AA06AB4CB77BBA7CDC6BCEE53C020B3343B9BD9A8298AD2055EE1A6070849140A86288721815C79734773F4097CF4741CC9635A30C8100B20733D3980B350393FAAC4CD0E66E4737C681DBBCC8D7953FA77454C422AD870E278B1121C33C8273370E5B686A6AAB17FCA3B67A3040D6491241BF5E3072FBDC1E422413FA5B4E9EE91EB3C936E21A5C7856942F44A55670A688A69E91A9A80BF4094C301DF705334DACB0CD929473829F34F37947D22B55C062F4CCF703EE3C1CC0BA7316DD658E6B6E0815F8FC9A70B1BBA325EC32E293091688A8FD05CD6DA066D2BAB105299B3EE66605BD5A803760AF56A6033CB9D3B9240A064D6C06CEAB73E59CFCA9FF6402255A326AEF1E9CB678BF36929DAFE29A58";

    // Iterate through KATs and validate
    foreach (keygen_kats[i]) begin
      parse_hex_to_array(keygen_kats[i].seed_d, kat_seed_d);
      parse_hex_to_array(keygen_kats[i].seed_z, kat_seed_z);
      parse_hex_to_array(keygen_kats[i].expected_PK, PK);
      parse_hex_to_array(keygen_kats[i].expected_SK, SK);

      `uvm_info("KAT", $sformatf("Running KeyGen KAT %0d", i), UVM_LOW);

      // Wait for ready flag in MLKEM_STATUS
      ready = 0;
      while (!ready) begin
        reg_model.MLKEM_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", "Failed to read MLKEM_STATUS");
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("MLKEM_STATUS: %h", data), UVM_HIGH);
        end
        ready = data[0];
      end

      // Write SEED to ML_KEM_SEED_D registers
      foreach (reg_model.MLKEM_SEED_D[j]) begin
        reg_model.MLKEM_SEED_D[j].write(status, kat_seed_d[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLKEM_SEED_D[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLKEM_SEED_D[%0d]: %h", j, kat_seed_d[j]), UVM_LOW);
        end
      end

      // Write SEED to ML_KEM_SEED_Z registers
      foreach (reg_model.MLKEM_SEED_Z[j]) begin
        reg_model.MLKEM_SEED_Z[j].write(status, kat_seed_z[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLKEM_SEED_Z[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLKEM_SEED_Z[%0d]: %h", j, kat_seed_z[j]), UVM_LOW);
        end
      end

      // Trigger KeyGen operation
      data = 'h00000001; // KeyGen command
      reg_model.MLKEM_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE_FAIL", "Failed to write MLKEM_CTRL to trigger KeyGen");
      end else begin
        `uvm_info("REG_WRITE_PASS", "Successfully wrote MLKEM_CTRL to trigger KeyGen", UVM_LOW);
      end

      // Wait for ready flag in MLKEM_STATUS
      valid =0;
      while(!valid) begin
        reg_model.MLKEM_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end
/*
      // Reading MLKEM_ENCAPS_KEY register
      for(int i = 0; i < reg_model.MLKEM_ENCAPS_KEY.m_mem.get_size(); i++) begin
        reg_model.MLKEM_ENCAPS_KEY.m_mem.read(status, i, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_ENCAPS_KEY[%0d]", i));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_ENCAPS_KEY[%0d]: %0h", i, data), UVM_LOW);
          if (PK[i] != data)
          `uvm_error("REG_READ", $sformatf("MLKEM_ENCAPS_KEY[%0d] mismatch: actual=0x%08h, expected=0x%08h",
                    i, data, PK[i]));
        end
      end
*/
      // Reading MLKEM_DECAPS_KEY register
      for(int i = 0; i < reg_model.MLKEM_DECAPS_KEY.m_mem.get_size(); i++) begin
        reg_model.MLKEM_DECAPS_KEY.m_mem.read(status, i, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_DECAPS_KEY[%0d]", i));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_DECAPS_KEY[%0d]: %0h", i, data), UVM_LOW);
          if (SK[i] != data)
          `uvm_error("REG_READ", $sformatf("MLKEM_DECAPS_KEY[%0d] mismatch: actual=0x%08h, expected=0x%08h",
                    i, data, SK[i]));
        end
      end

      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end

    `uvm_info("KAT", $sformatf("KeyGen KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



