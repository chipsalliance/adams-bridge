
// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
import uvm_pkg::*;

`uvm_analysis_imp_decl(_ntt_txn)
`uvm_analysis_imp_decl(_ntt_mem_txn)
`uvm_analysis_imp_decl(_pwm_a_mem_txn)
`uvm_analysis_imp_decl(_pwm_b_mem_txn)

parameter logic [22:0] zetas[0:255] = '{
    23'd1,
    23'd4808194,
    23'd3765607,
    23'd3761513,
    23'd5178923,
    23'd5496691,
    23'd5234739,
    23'd5178987,
    23'd7778734,
    23'd3542485,
    23'd2682288,
    23'd2129892,
    23'd3764867,
    23'd7375178,
    23'd557458,
    23'd7159240,
    23'd5010068,
    23'd4317364,
    23'd2663378,
    23'd6705802,
    23'd4855975,
    23'd7946292,
    23'd676590,
    23'd7044481,
    23'd5152541,
    23'd1714295,
    23'd2453983,
    23'd1460718,
    23'd7737789,
    23'd4795319,
    23'd2815639,
    23'd2283733,
    23'd3602218,
    23'd3182878,
    23'd2740543,
    23'd4793971,
    23'd5269599,
    23'd2101410,
    23'd3704823,
    23'd1159875,
    23'd394148,
    23'd928749,
    23'd1095468,
    23'd4874037,
    23'd2071829,
    23'd4361428,
    23'd3241972,
    23'd2156050,
    23'd3415069,
    23'd1759347,
    23'd7562881,
    23'd4805951,
    23'd3756790,
    23'd6444618,
    23'd6663429,
    23'd4430364,
    23'd5483103,
    23'd3192354,
    23'd556856,
    23'd3870317,
    23'd2917338,
    23'd1853806,
    23'd3345963,
    23'd1858416,
    23'd3073009,
    23'd1277625,
    23'd5744944,
    23'd3852015,
    23'd4183372,
    23'd5157610,
    23'd5258977,
    23'd8106357,
    23'd2508980,
    23'd2028118,
    23'd1937570,
    23'd4564692,
    23'd2811291,
    23'd5396636,
    23'd7270901,
    23'd4158088,
    23'd1528066,
    23'd482649,
    23'd1148858,
    23'd5418153,
    23'd7814814,
    23'd169688,
    23'd2462444,
    23'd5046034,
    23'd4213992,
    23'd4892034,
    23'd1987814,
    23'd5183169,
    23'd1736313,
    23'd235407,
    23'd5130263,
    23'd3258457,
    23'd5801164,
    23'd1787943,
    23'd5989328,
    23'd6125690,
    23'd3482206,
    23'd4197502,
    23'd7080401,
    23'd6018354,
    23'd7062739,
    23'd2461387,
    23'd3035980,
    23'd621164,
    23'd3901472,
    23'd7153756,
    23'd2925816,
    23'd3374250,
    23'd1356448,
    23'd5604662,
    23'd2683270,
    23'd5601629,
    23'd4912752,
    23'd2312838,
    23'd7727142,
    23'd7921254,
    23'd348812,
    23'd8052569,
    23'd1011223,
    23'd6026202,
    23'd4561790,
    23'd6458164,
    23'd6143691,
    23'd1744507,
    23'd1753,
    23'd6444997,
    23'd5720892,
    23'd6924527,
    23'd2660408,
    23'd6600190,
    23'd8321269,
    23'd2772600,
    23'd1182243,
    23'd87208,
    23'd636927,
    23'd4415111,
    23'd4423672,
    23'd6084020,
    23'd5095502,
    23'd4663471,
    23'd8352605,
    23'd822541,
    23'd1009365,
    23'd5926272,
    23'd6400920,
    23'd1596822,
    23'd4423473,
    23'd4620952,
    23'd6695264,
    23'd4969849,
    23'd2678278,
    23'd4611469,
    23'd4829411,
    23'd635956,
    23'd8129971,
    23'd5925040,
    23'd4234153,
    23'd6607829,
    23'd2192938,
    23'd6653329,
    23'd2387513,
    23'd4768667,
    23'd8111961,
    23'd5199961,
    23'd3747250,
    23'd2296099,
    23'd1239911,
    23'd4541938,
    23'd3195676,
    23'd2642980,
    23'd1254190,
    23'd8368000,
    23'd2998219,
    23'd141835,
    23'd8291116,
    23'd2513018,
    23'd7025525,
    23'd613238,
    23'd7070156,
    23'd6161950,
    23'd7921677,
    23'd6458423,
    23'd4040196,
    23'd4908348,
    23'd2039144,
    23'd6500539,
    23'd7561656,
    23'd6201452,
    23'd6757063,
    23'd2105286,
    23'd6006015,
    23'd6346610,
    23'd586241,
    23'd7200804,
    23'd527981,
    23'd5637006,
    23'd6903432,
    23'd1994046,
    23'd2491325,
    23'd6987258,
    23'd507927,
    23'd7192532,
    23'd7655613,
    23'd6545891,
    23'd5346675,
    23'd8041997,
    23'd2647994,
    23'd3009748,
    23'd5767564,
    23'd4148469,
    23'd749577,
    23'd4357667,
    23'd3980599,
    23'd2569011,
    23'd6764887,
    23'd1723229,
    23'd1665318,
    23'd2028038,
    23'd1163598,
    23'd5011144,
    23'd3994671,
    23'd8368538,
    23'd7009900,
    23'd3020393,
    23'd3363542,
    23'd214880,
    23'd545376,
    23'd7609976,
    23'd3105558,
    23'd7277073,
    23'd508145,
    23'd7826699,
    23'd860144,
    23'd3430436,
    23'd140244,
    23'd6866265,
    23'd6195333,
    23'd3123762,
    23'd2358373,
    23'd6187330,
    23'd5365997,
    23'd6663603,
    23'd2926054,
    23'd7987710,
    23'd8077412,
    23'd3531229,
    23'd4405932,
    23'd4606686,
    23'd1900052,
    23'd7598542,
    23'd1054478,
    23'd7648983
};

logic [23:0] zetas_inv[0:255] = '{
    23'd8380416,
    23'd3572223,
    23'd4614810,
    23'd4618904,
    23'd3201494,
    23'd2883726,
    23'd3145678,
    23'd3201430,
    23'd601683,
    23'd4837932,
    23'd5698129,
    23'd6250525,
    23'd4615550,
    23'd1005239,
    23'd7822959,
    23'd1221177,
    23'd3370349,
    23'd4063053,
    23'd5717039,
    23'd1674615,
    23'd3524442,
    23'd434125,
    23'd7703827,
    23'd1335936,
    23'd3227876,
    23'd6666122,
    23'd5926434,
    23'd6919699,
    23'd642628,
    23'd3585098,
    23'd5564778,
    23'd6096684,
    23'd4778199,
    23'd5197539,
    23'd5639874,
    23'd3586446,
    23'd3110818,
    23'd6279007,
    23'd4675594,
    23'd7220542,
    23'd7986269,
    23'd7451668,
    23'd7284949,
    23'd3506380,
    23'd6308588,
    23'd4018989,
    23'd5138445,
    23'd6224367,
    23'd4965348,
    23'd6621070,
    23'd817536,
    23'd3574466,
    23'd4623627,
    23'd1935799,
    23'd1716988,
    23'd3950053,
    23'd2897314,
    23'd5188063,
    23'd7823561,
    23'd4510100,
    23'd5463079,
    23'd6526611,
    23'd5034454,
    23'd6522001,
    23'd5307408,
    23'd7102792,
    23'd2635473,
    23'd4528402,
    23'd4197045,
    23'd3222807,
    23'd3121440,
    23'd274060,
    23'd5871437,
    23'd6352299,
    23'd6442847,
    23'd3815725,
    23'd5569126,
    23'd2983781,
    23'd1109516,
    23'd4222329,
    23'd6852351,
    23'd7897768,
    23'd7231559,
    23'd2962264,
    23'd565603,
    23'd8210729,
    23'd5917973,
    23'd3334383,
    23'd4166425,
    23'd3488383,
    23'd6392603,
    23'd3197248,
    23'd6644104,
    23'd8145010,
    23'd3250154,
    23'd5121960,
    23'd2579253,
    23'd6592474,
    23'd2391089,
    23'd2254727,
    23'd4898211,
    23'd4182915,
    23'd1300016,
    23'd2362063,
    23'd1317678,
    23'd5919030,
    23'd5344437,
    23'd7759253,
    23'd4478945,
    23'd1226661,
    23'd5454601,
    23'd5006167,
    23'd7023969,
    23'd2775755,
    23'd5697147,
    23'd2778788,
    23'd3467665,
    23'd6067579,
    23'd653275,
    23'd459163,
    23'd8031605,
    23'd327848,
    23'd7369194,
    23'd2354215,
    23'd3818627,
    23'd1922253,
    23'd2236726,
    23'd6635910,
    23'd8378664,
    23'd1935420,
    23'd2659525,
    23'd1455890,
    23'd5720009,
    23'd1780227,
    23'd59148,
    23'd5607817,
    23'd7198174,
    23'd8293209,
    23'd7743490,
    23'd3965306,
    23'd3956745,
    23'd2296397,
    23'd3284915,
    23'd3716946,
    23'd27812,
    23'd7557876,
    23'd7371052,
    23'd2454145,
    23'd1979497,
    23'd6783595,
    23'd3956944,
    23'd3759465,
    23'd1685153,
    23'd3410568,
    23'd5702139,
    23'd3768948,
    23'd3551006,
    23'd7744461,
    23'd250446,
    23'd2455377,
    23'd4146264,
    23'd1772588,
    23'd6187479,
    23'd1727088,
    23'd5992904,
    23'd3611750,
    23'd268456,
    23'd3180456,
    23'd4633167,
    23'd6084318,
    23'd7140506,
    23'd3838479,
    23'd5184741,
    23'd5737437,
    23'd7126227,
    23'd12417,
    23'd5382198,
    23'd8238582,
    23'd89301,
    23'd5867399,
    23'd1354892,
    23'd7767179,
    23'd1310261,
    23'd2218467,
    23'd458740,
    23'd1921994,
    23'd4340221,
    23'd3472069,
    23'd6341273,
    23'd1879878,
    23'd818761,
    23'd2178965,
    23'd1623354,
    23'd6275131,
    23'd2374402,
    23'd2033807,
    23'd7794176,
    23'd1179613,
    23'd7852436,
    23'd2743411,
    23'd1476985,
    23'd6386371,
    23'd5889092,
    23'd1393159,
    23'd7872490,
    23'd1187885,
    23'd724804,
    23'd1834526,
    23'd3033742,
    23'd338420,
    23'd5732423,
    23'd5370669,
    23'd2612853,
    23'd4231948,
    23'd7630840,
    23'd4022750,
    23'd4399818,
    23'd5811406,
    23'd1615530,
    23'd6657188,
    23'd6715099,
    23'd6352379,
    23'd7216819,
    23'd3369273,
    23'd4385746,
    23'd11879,
    23'd1370517,
    23'd5360024,
    23'd5016875,
    23'd8165537,
    23'd7835041,
    23'd770441,
    23'd5274859,
    23'd1103344,
    23'd7872272,
    23'd553718,
    23'd7520273,
    23'd4949981,
    23'd8240173,
    23'd1514152,
    23'd2185084,
    23'd5256655,
    23'd6022044,
    23'd2193087,
    23'd3014420,
    23'd1716814,
    23'd5454363,
    23'd392707,
    23'd303005,
    23'd4849188,
    23'd3974485,
    23'd3773731,
    23'd6480365,
    23'd781875,
    23'd7325939,
    23'd731434
};