// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
//======================================================================
//
// twiddle_rom.sv
// --------
// ROM contains twiddle factors for NTT and INTT
// 
//
//======================================================================

module ntt_twiddle_lookup 
    import ntt_defines_pkg::*;
#(
    parameter ADDR_WIDTH = 7,
    parameter DATA_WIDTH = 24,
    parameter KYBER_DATA_WIDTH = 12
)
(

    input mode_t mode,
    input wire [ADDR_WIDTH-1:0] raddr,
    input wire mlkem,
    output logic [(3*DATA_WIDTH)-1:0] rdata
);

reg [(3*DATA_WIDTH)-1:0] ntt_twiddle_mem  [84:0];
reg [(3*DATA_WIDTH)-1:0] intt_twiddle_mem [84:0];
reg [(3*KYBER_DATA_WIDTH)-1:0] kyber_ntt_twiddle_mem  [84:0];
reg [(3*KYBER_DATA_WIDTH)-1:0] kyber_intt_twiddle_mem [84:0];

always_comb begin
    if (mlkem) //TODO: make sure there is no pairwm op after gs
        rdata = (mode inside {ct, pwm}) ? {12'h0, kyber_ntt_twiddle_mem[raddr]} : (mode == gs) ? {12'h0, kyber_intt_twiddle_mem[raddr]} : 'h0;
    else
        rdata = (mode == ct) ? ntt_twiddle_mem[raddr] : (mode == gs) ? intt_twiddle_mem[raddr] : 'h0;
end

logic [255 : 0][(DATA_WIDTH)-1:0] zeta;
logic [255 : 0][(DATA_WIDTH)-1:0] zetainv;
logic [255 : 0][KYBER_DATA_WIDTH-1:0] kyber_zeta;
logic [255 : 0][KYBER_DATA_WIDTH-1:0] kyber_zetainv;

assign zeta[0] = 23'h000001;
assign zeta[1] = 23'h495E02;
assign zeta[2] = 23'h397567;
assign zeta[3] = 23'h396569;
assign zeta[4] = 23'h4F062B;
assign zeta[5] = 23'h53DF73;
assign zeta[6] = 23'h4FE033;
assign zeta[7] = 23'h4F066B;
assign zeta[8] = 23'h76B1AE;
assign zeta[9] = 23'h360DD5;
assign zeta[10] = 23'h28EDB0;
assign zeta[11] = 23'h207FE4;
assign zeta[12] = 23'h397283;
assign zeta[13] = 23'h70894A;
assign zeta[14] = 23'h088192;
assign zeta[15] = 23'h6D3DC8;
assign zeta[16] = 23'h4C7294;
assign zeta[17] = 23'h41E0B4;
assign zeta[18] = 23'h28A3D2;
assign zeta[19] = 23'h66528A;
assign zeta[20] = 23'h4A18A7;
assign zeta[21] = 23'h794034;
assign zeta[22] = 23'h0A52EE;
assign zeta[23] = 23'h6B7D81;
assign zeta[24] = 23'h4E9F1D;
assign zeta[25] = 23'h1A2877;
assign zeta[26] = 23'h2571DF;
assign zeta[27] = 23'h1649EE;
assign zeta[28] = 23'h7611BD;
assign zeta[29] = 23'h492BB7;
assign zeta[30] = 23'h2AF697;
assign zeta[31] = 23'h22D8D5;
assign zeta[32] = 23'h36F72A;
assign zeta[33] = 23'h30911E;
assign zeta[34] = 23'h29D13F;
assign zeta[35] = 23'h492673;
assign zeta[36] = 23'h50685F;
assign zeta[37] = 23'h2010A2;
assign zeta[38] = 23'h3887F7;
assign zeta[39] = 23'h11B2C3;
assign zeta[40] = 23'h0603A4;
assign zeta[41] = 23'h0E2BED;
assign zeta[42] = 23'h10B72C;
assign zeta[43] = 23'h4A5F35;
assign zeta[44] = 23'h1F9D15;
assign zeta[45] = 23'h428CD4;
assign zeta[46] = 23'h3177F4;
assign zeta[47] = 23'h20E612;
assign zeta[48] = 23'h341C1D;
assign zeta[49] = 23'h1AD873;
assign zeta[50] = 23'h736681;
assign zeta[51] = 23'h49553F;
assign zeta[52] = 23'h3952F6;
assign zeta[53] = 23'h62564A;
assign zeta[54] = 23'h65AD05;
assign zeta[55] = 23'h439A1C;
assign zeta[56] = 23'h53AA5F;
assign zeta[57] = 23'h30B622;
assign zeta[58] = 23'h087F38;
assign zeta[59] = 23'h3B0E6D;
assign zeta[60] = 23'h2C83DA;
assign zeta[61] = 23'h1C496E;
assign zeta[62] = 23'h330E2B;
assign zeta[63] = 23'h1C5B70;
assign zeta[64] = 23'h2EE3F1;
assign zeta[65] = 23'h137EB9;
assign zeta[66] = 23'h57A930;
assign zeta[67] = 23'h3AC6EF;
assign zeta[68] = 23'h3FD54C;
assign zeta[69] = 23'h4EB2EA;
assign zeta[70] = 23'h503EE1;
assign zeta[71] = 23'h7BB175;
assign zeta[72] = 23'h2648B4;
assign zeta[73] = 23'h1EF256;
assign zeta[74] = 23'h1D90A2;
assign zeta[75] = 23'h45A6D4;
assign zeta[76] = 23'h2AE59B;
assign zeta[77] = 23'h52589C;
assign zeta[78] = 23'h6EF1F5;
assign zeta[79] = 23'h3F7288;
assign zeta[80] = 23'h175102;
assign zeta[81] = 23'h075D59;
assign zeta[82] = 23'h1187BA;
assign zeta[83] = 23'h52ACA9;
assign zeta[84] = 23'h773E9E;
assign zeta[85] = 23'h0296D8;
assign zeta[86] = 23'h2592EC;
assign zeta[87] = 23'h4CFF12;
assign zeta[88] = 23'h404CE8;
assign zeta[89] = 23'h4AA582;
assign zeta[90] = 23'h1E54E6;
assign zeta[91] = 23'h4F16C1;
assign zeta[92] = 23'h1A7E79;
assign zeta[93] = 23'h03978F;
assign zeta[94] = 23'h4E4817;
assign zeta[95] = 23'h31B859;
assign zeta[96] = 23'h5884CC;
assign zeta[97] = 23'h1B4827;
assign zeta[98] = 23'h5B63D0;
assign zeta[99] = 23'h5D787A;
assign zeta[100] = 23'h35225E;
assign zeta[101] = 23'h400C7E;
assign zeta[102] = 23'h6C09D1;
assign zeta[103] = 23'h5BD532;
assign zeta[104] = 23'h6BC4D3;
assign zeta[105] = 23'h258ECB;
assign zeta[106] = 23'h2E534C;
assign zeta[107] = 23'h097A6C;
assign zeta[108] = 23'h3B8820;
assign zeta[109] = 23'h6D285C;
assign zeta[110] = 23'h2CA4F8;
assign zeta[111] = 23'h337CAA;
assign zeta[112] = 23'h14B2A0;
assign zeta[113] = 23'h558536;
assign zeta[114] = 23'h28F186;
assign zeta[115] = 23'h55795D;
assign zeta[116] = 23'h4AF670;
assign zeta[117] = 23'h234A86;
assign zeta[118] = 23'h75E826;
assign zeta[119] = 23'h78DE66;
assign zeta[120] = 23'h05528C;
assign zeta[121] = 23'h7ADF59;
assign zeta[122] = 23'h0F6E17;
assign zeta[123] = 23'h5BF3DA;
assign zeta[124] = 23'h459B7E;
assign zeta[125] = 23'h628B34;
assign zeta[126] = 23'h5DBECB;
assign zeta[127] = 23'h1A9E7B;
assign zeta[128] = 23'h0006D9;
assign zeta[129] = 23'h6257C5;
assign zeta[130] = 23'h574B3C;
assign zeta[131] = 23'h69A8EF;
assign zeta[132] = 23'h289838;
assign zeta[133] = 23'h64B5FE;
assign zeta[134] = 23'h7EF8F5;
assign zeta[135] = 23'h2A4E78;
assign zeta[136] = 23'h120A23;
assign zeta[137] = 23'h0154A8;
assign zeta[138] = 23'h09B7FF;
assign zeta[139] = 23'h435E87;
assign zeta[140] = 23'h437FF8;
assign zeta[141] = 23'h5CD5B4;
assign zeta[142] = 23'h4DC04E;
assign zeta[143] = 23'h4728AF;
assign zeta[144] = 23'h7F735D;
assign zeta[145] = 23'h0C8D0D;
assign zeta[146] = 23'h0F66D5;
assign zeta[147] = 23'h5A6D80;
assign zeta[148] = 23'h61AB98;
assign zeta[149] = 23'h185D96;
assign zeta[150] = 23'h437F31;
assign zeta[151] = 23'h468298;
assign zeta[152] = 23'h662960;
assign zeta[153] = 23'h4BD579;
assign zeta[154] = 23'h28DE06;
assign zeta[155] = 23'h465D8D;
assign zeta[156] = 23'h49B0E3;
assign zeta[157] = 23'h09B434;
assign zeta[158] = 23'h7C0DB3;
assign zeta[159] = 23'h5A68B0;
assign zeta[160] = 23'h409BA9;
assign zeta[161] = 23'h64D3D5;
assign zeta[162] = 23'h21762A;
assign zeta[163] = 23'h658591;
assign zeta[164] = 23'h246E39;
assign zeta[165] = 23'h48C39B;
assign zeta[166] = 23'h7BC759;
assign zeta[167] = 23'h4F5859;
assign zeta[168] = 23'h392DB2;
assign zeta[169] = 23'h230923;
assign zeta[170] = 23'h12EB67;
assign zeta[171] = 23'h454DF2;
assign zeta[172] = 23'h30C31C;
assign zeta[173] = 23'h285424;
assign zeta[174] = 23'h13232E;
assign zeta[175] = 23'h7FAF80;
assign zeta[176] = 23'h2DBFCB;
assign zeta[177] = 23'h022A0B;
assign zeta[178] = 23'h7E832C;
assign zeta[179] = 23'h26587A;
assign zeta[180] = 23'h6B3375;
assign zeta[181] = 23'h095B76;
assign zeta[182] = 23'h6BE1CC;
assign zeta[183] = 23'h5E061E;
assign zeta[184] = 23'h78E00D;
assign zeta[185] = 23'h628C37;
assign zeta[186] = 23'h3DA604;
assign zeta[187] = 23'h4AE53C;
assign zeta[188] = 23'h1F1D68;
assign zeta[189] = 23'h6330BB;
assign zeta[190] = 23'h7361B8;
assign zeta[191] = 23'h5EA06C;
assign zeta[192] = 23'h671AC7;
assign zeta[193] = 23'h201FC6;
assign zeta[194] = 23'h5BA4FF;
assign zeta[195] = 23'h60D772;
assign zeta[196] = 23'h08F201;
assign zeta[197] = 23'h6DE024;
assign zeta[198] = 23'h080E6D;
assign zeta[199] = 23'h56038E;
assign zeta[200] = 23'h695688;
assign zeta[201] = 23'h1E6D3E;
assign zeta[202] = 23'h2603BD;
assign zeta[203] = 23'h6A9DFA;
assign zeta[204] = 23'h07C017;
assign zeta[205] = 23'h6DBFD4;
assign zeta[206] = 23'h74D0BD;
assign zeta[207] = 23'h63E1E3;
assign zeta[208] = 23'h519573;
assign zeta[209] = 23'h7AB60D;
assign zeta[210] = 23'h2867BA;
assign zeta[211] = 23'h2DECD4;
assign zeta[212] = 23'h58018C;
assign zeta[213] = 23'h3F4CF5;
assign zeta[214] = 23'h0B7009;
assign zeta[215] = 23'h427E23;
assign zeta[216] = 23'h3CBD37;
assign zeta[217] = 23'h273333;
assign zeta[218] = 23'h673957;
assign zeta[219] = 23'h1A4B5D;
assign zeta[220] = 23'h196926;
assign zeta[221] = 23'h1EF206;
assign zeta[222] = 23'h11C14E;
assign zeta[223] = 23'h4C76C8;
assign zeta[224] = 23'h3CF42F;
assign zeta[225] = 23'h7FB19A;
assign zeta[226] = 23'h6AF66C;
assign zeta[227] = 23'h2E1669;
assign zeta[228] = 23'h3352D6;
assign zeta[229] = 23'h034760;
assign zeta[230] = 23'h085260;
assign zeta[231] = 23'h741E78;
assign zeta[232] = 23'h2F6316;
assign zeta[233] = 23'h6F0A11;
assign zeta[234] = 23'h07C0F1;
assign zeta[235] = 23'h776D0B;
assign zeta[236] = 23'h0D1FF0;
assign zeta[237] = 23'h345824;
assign zeta[238] = 23'h0223D4;
assign zeta[239] = 23'h68C559;
assign zeta[240] = 23'h5E8885;
assign zeta[241] = 23'h2FAA32;
assign zeta[242] = 23'h23FC65;
assign zeta[243] = 23'h5E6942;
assign zeta[244] = 23'h51E0ED;
assign zeta[245] = 23'h65ADB3;
assign zeta[246] = 23'h2CA5E6;
assign zeta[247] = 23'h79E1FE;
assign zeta[248] = 23'h7B4064;
assign zeta[249] = 23'h35E1DD;
assign zeta[250] = 23'h433AAC;
assign zeta[251] = 23'h464ADE;
assign zeta[252] = 23'h1CFE14;
assign zeta[253] = 23'h73F1CE;
assign zeta[254] = 23'h10170E;
assign zeta[255] = 23'h74B6D7;

//------------------------------------------------------------------------------------


assign zetainv[0] = 23'h7FE000;
assign zetainv[1] = 23'h3681FF;
assign zetainv[2] = 23'h466A9A;
assign zetainv[3] = 23'h467A98;
assign zetainv[4] = 23'h30D9D6;
assign zetainv[5] = 23'h2C008E;
assign zetainv[6] = 23'h2FFFCE;
assign zetainv[7] = 23'h30D996;
assign zetainv[8] = 23'h092E53;
assign zetainv[9] = 23'h49D22C;
assign zetainv[10] = 23'h56F251;
assign zetainv[11] = 23'h5F601D;
assign zetainv[12] = 23'h466D7E;
assign zetainv[13] = 23'h0F56B7;
assign zetainv[14] = 23'h775E6F;
assign zetainv[15] = 23'h12A239;
assign zetainv[16] = 23'h336D6D;
assign zetainv[17] = 23'h3DFF4D;
assign zetainv[18] = 23'h573C2F;
assign zetainv[19] = 23'h198D77;
assign zetainv[20] = 23'h35C75A;
assign zetainv[21] = 23'h069FCD;
assign zetainv[22] = 23'h758D13;
assign zetainv[23] = 23'h146280;
assign zetainv[24] = 23'h3140E4;
assign zetainv[25] = 23'h65B78A;
assign zetainv[26] = 23'h5A6E22;
assign zetainv[27] = 23'h699613;
assign zetainv[28] = 23'h09CE44;
assign zetainv[29] = 23'h36B44A;
assign zetainv[30] = 23'h54E96A;
assign zetainv[31] = 23'h5D072C;
assign zetainv[32] = 23'h48E8D7;
assign zetainv[33] = 23'h4F4EE3;
assign zetainv[34] = 23'h560EC2;
assign zetainv[35] = 23'h36B98E;
assign zetainv[36] = 23'h2F77A2;
assign zetainv[37] = 23'h5FCF5F;
assign zetainv[38] = 23'h47580A;
assign zetainv[39] = 23'h6E2D3E;
assign zetainv[40] = 23'h79DC5D;
assign zetainv[41] = 23'h71B414;
assign zetainv[42] = 23'h6F28D5;
assign zetainv[43] = 23'h3580CC;
assign zetainv[44] = 23'h6042EC;
assign zetainv[45] = 23'h3D532D;
assign zetainv[46] = 23'h4E680D;
assign zetainv[47] = 23'h5EF9EF;
assign zetainv[48] = 23'h4BC3E4;
assign zetainv[49] = 23'h65078E;
assign zetainv[50] = 23'h0C7980;
assign zetainv[51] = 23'h368AC2;
assign zetainv[52] = 23'h468D0B;
assign zetainv[53] = 23'h1D89B7;
assign zetainv[54] = 23'h1A32FC;
assign zetainv[55] = 23'h3C45E5;
assign zetainv[56] = 23'h2C35A2;
assign zetainv[57] = 23'h4F29DF;
assign zetainv[58] = 23'h7760C9;
assign zetainv[59] = 23'h44D194;
assign zetainv[60] = 23'h535C27;
assign zetainv[61] = 23'h639693;
assign zetainv[62] = 23'h4CD1D6;
assign zetainv[63] = 23'h638491;
assign zetainv[64] = 23'h50FC10;
assign zetainv[65] = 23'h6C6148;
assign zetainv[66] = 23'h2836D1;
assign zetainv[67] = 23'h451912;
assign zetainv[68] = 23'h400AB5;
assign zetainv[69] = 23'h312D17;
assign zetainv[70] = 23'h2FA120;
assign zetainv[71] = 23'h042E8C;
assign zetainv[72] = 23'h59974D;
assign zetainv[73] = 23'h60EDAB;
assign zetainv[74] = 23'h624F5F;
assign zetainv[75] = 23'h3A392D;
assign zetainv[76] = 23'h54FA66;
assign zetainv[77] = 23'h2D8765;
assign zetainv[78] = 23'h10EE0C;
assign zetainv[79] = 23'h406D79;
assign zetainv[80] = 23'h688EFF;
assign zetainv[81] = 23'h7882A8;
assign zetainv[82] = 23'h6E5847;
assign zetainv[83] = 23'h2D3358;
assign zetainv[84] = 23'h08A163;
assign zetainv[85] = 23'h7D4929;
assign zetainv[86] = 23'h5A4D15;
assign zetainv[87] = 23'h32E0EF;
assign zetainv[88] = 23'h3F9319;
assign zetainv[89] = 23'h353A7F;
assign zetainv[90] = 23'h618B1B;
assign zetainv[91] = 23'h30C940;
assign zetainv[92] = 23'h656188;
assign zetainv[93] = 23'h7C4872;
assign zetainv[94] = 23'h3197EA;
assign zetainv[95] = 23'h4E27A8;
assign zetainv[96] = 23'h275B35;
assign zetainv[97] = 23'h6497DA;
assign zetainv[98] = 23'h247C31;
assign zetainv[99] = 23'h226787;
assign zetainv[100] = 23'h4ABDA3;
assign zetainv[101] = 23'h3FD383;
assign zetainv[102] = 23'h13D630;
assign zetainv[103] = 23'h240ACF;
assign zetainv[104] = 23'h141B2E;
assign zetainv[105] = 23'h5A5136;
assign zetainv[106] = 23'h518CB5;
assign zetainv[107] = 23'h766595;
assign zetainv[108] = 23'h4457E1;
assign zetainv[109] = 23'h12B7A5;
assign zetainv[110] = 23'h533B09;
assign zetainv[111] = 23'h4C6357;
assign zetainv[112] = 23'h6B2D61;
assign zetainv[113] = 23'h2A5ACB;
assign zetainv[114] = 23'h56EE7B;
assign zetainv[115] = 23'h2A66A4;
assign zetainv[116] = 23'h34E991;
assign zetainv[117] = 23'h5C957B;
assign zetainv[118] = 23'h09F7DB;
assign zetainv[119] = 23'h07019B;
assign zetainv[120] = 23'h7A8D75;
assign zetainv[121] = 23'h0500A8;
assign zetainv[122] = 23'h7071EA;
assign zetainv[123] = 23'h23EC27;
assign zetainv[124] = 23'h3A4483;
assign zetainv[125] = 23'h1D54CD;
assign zetainv[126] = 23'h222136;
assign zetainv[127] = 23'h654186;
assign zetainv[128] = 23'h7FD928;
assign zetainv[129] = 23'h1D883C;
assign zetainv[130] = 23'h2894C5;
assign zetainv[131] = 23'h163712;
assign zetainv[132] = 23'h5747C9;
assign zetainv[133] = 23'h1B2A03;
assign zetainv[134] = 23'h00E70C;
assign zetainv[135] = 23'h559189;
assign zetainv[136] = 23'h6DD5DE;
assign zetainv[137] = 23'h7E8B59;
assign zetainv[138] = 23'h762802;
assign zetainv[139] = 23'h3C817A;
assign zetainv[140] = 23'h3C6009;
assign zetainv[141] = 23'h230A4D;
assign zetainv[142] = 23'h321FB3;
assign zetainv[143] = 23'h38B752;
assign zetainv[144] = 23'h006CA4;
assign zetainv[145] = 23'h7352F4;
assign zetainv[146] = 23'h70792C;
assign zetainv[147] = 23'h257281;
assign zetainv[148] = 23'h1E3469;
assign zetainv[149] = 23'h67826B;
assign zetainv[150] = 23'h3C60D0;
assign zetainv[151] = 23'h395D69;
assign zetainv[152] = 23'h19B6A1;
assign zetainv[153] = 23'h340A88;
assign zetainv[154] = 23'h5701FB;
assign zetainv[155] = 23'h398274;
assign zetainv[156] = 23'h362F1E;
assign zetainv[157] = 23'h762BCD;
assign zetainv[158] = 23'h03D24E;
assign zetainv[159] = 23'h257751;
assign zetainv[160] = 23'h3F4458;
assign zetainv[161] = 23'h1B0C2C;
assign zetainv[162] = 23'h5E69D7;
assign zetainv[163] = 23'h1A5A70;
assign zetainv[164] = 23'h5B71C8;
assign zetainv[165] = 23'h371C66;
assign zetainv[166] = 23'h0418A8;
assign zetainv[167] = 23'h3087A8;
assign zetainv[168] = 23'h46B24F;
assign zetainv[169] = 23'h5CD6DE;
assign zetainv[170] = 23'h6CF49A;
assign zetainv[171] = 23'h3A920F;
assign zetainv[172] = 23'h4F1CE5;
assign zetainv[173] = 23'h578BDD;
assign zetainv[174] = 23'h6CBCD3;
assign zetainv[175] = 23'h003081;
assign zetainv[176] = 23'h522036;
assign zetainv[177] = 23'h7DB5F6;
assign zetainv[178] = 23'h015CD5;
assign zetainv[179] = 23'h598787;
assign zetainv[180] = 23'h14AC8C;
assign zetainv[181] = 23'h76848B;
assign zetainv[182] = 23'h13FE35;
assign zetainv[183] = 23'h21D9E3;
assign zetainv[184] = 23'h06FFF4;
assign zetainv[185] = 23'h1D53CA;
assign zetainv[186] = 23'h4239FD;
assign zetainv[187] = 23'h34FAC5;
assign zetainv[188] = 23'h60C299;
assign zetainv[189] = 23'h1CAF46;
assign zetainv[190] = 23'h0C7E49;
assign zetainv[191] = 23'h213F95;
assign zetainv[192] = 23'h18C53A;
assign zetainv[193] = 23'h5FC03B;
assign zetainv[194] = 23'h243B02;
assign zetainv[195] = 23'h1F088F;
assign zetainv[196] = 23'h76EE00;
assign zetainv[197] = 23'h11FFDD;
assign zetainv[198] = 23'h77D194;
assign zetainv[199] = 23'h29DC73;
assign zetainv[200] = 23'h168979;
assign zetainv[201] = 23'h6172C3;
assign zetainv[202] = 23'h59DC44;
assign zetainv[203] = 23'h154207;
assign zetainv[204] = 23'h781FEA;
assign zetainv[205] = 23'h12202D;
assign zetainv[206] = 23'h0B0F44;
assign zetainv[207] = 23'h1BFE1E;
assign zetainv[208] = 23'h2E4A8E;
assign zetainv[209] = 23'h0529F4;
assign zetainv[210] = 23'h577847;
assign zetainv[211] = 23'h51F32D;
assign zetainv[212] = 23'h27DE75;
assign zetainv[213] = 23'h40930C;
assign zetainv[214] = 23'h746FF8;
assign zetainv[215] = 23'h3D61DE;
assign zetainv[216] = 23'h4322CA;
assign zetainv[217] = 23'h58ACCE;
assign zetainv[218] = 23'h18A6AA;
assign zetainv[219] = 23'h6594A4;
assign zetainv[220] = 23'h6676DB;
assign zetainv[221] = 23'h60EDFB;
assign zetainv[222] = 23'h6E1EB3;
assign zetainv[223] = 23'h336939;
assign zetainv[224] = 23'h42EBD2;
assign zetainv[225] = 23'h002E67;
assign zetainv[226] = 23'h14E995;
assign zetainv[227] = 23'h51C998;
assign zetainv[228] = 23'h4C8D2B;
assign zetainv[229] = 23'h7C98A1;
assign zetainv[230] = 23'h778DA1;
assign zetainv[231] = 23'h0BC189;
assign zetainv[232] = 23'h507CEB;
assign zetainv[233] = 23'h10D5F0;
assign zetainv[234] = 23'h781F10;
assign zetainv[235] = 23'h0872F6;
assign zetainv[236] = 23'h72C011;
assign zetainv[237] = 23'h4B87DD;
assign zetainv[238] = 23'h7DBC2D;
assign zetainv[239] = 23'h171AA8;
assign zetainv[240] = 23'h21577C;
assign zetainv[241] = 23'h5035CF;
assign zetainv[242] = 23'h5BE39C;
assign zetainv[243] = 23'h2176BF;
assign zetainv[244] = 23'h2DFF14;
assign zetainv[245] = 23'h1A324E;
assign zetainv[246] = 23'h533A1B;
assign zetainv[247] = 23'h05FE03;
assign zetainv[248] = 23'h049F9D;
assign zetainv[249] = 23'h49FE24;
assign zetainv[250] = 23'h3CA555;
assign zetainv[251] = 23'h399523;
assign zetainv[252] = 23'h62E1ED;
assign zetainv[253] = 23'h0BEE33;
assign zetainv[254] = 23'h6FC8F3;
assign zetainv[255] = 23'h0B292A;

//------------------------------------------------------------------------------------

assign kyber_zeta[0]  = 12'h001 ;
assign kyber_zeta[1]  = 12'h6C1 ;
assign kyber_zeta[2]  = 12'hA14 ;
assign kyber_zeta[3]  = 12'hCD9 ;
assign kyber_zeta[4]  = 12'hA52 ;
assign kyber_zeta[5]  = 12'h276 ;
assign kyber_zeta[6]  = 12'h769 ;
assign kyber_zeta[7]  = 12'h350 ;
assign kyber_zeta[8]  = 12'h426 ;
assign kyber_zeta[9]  = 12'h77F ;
assign kyber_zeta[10] = 12'h0C1 ;
assign kyber_zeta[11] = 12'h31D ;
assign kyber_zeta[12] = 12'hAE2 ;
assign kyber_zeta[13] = 12'hCBC ;
assign kyber_zeta[14] = 12'h239 ;
assign kyber_zeta[15] = 12'h6D2 ;
assign kyber_zeta[16] = 12'h128 ;
assign kyber_zeta[17] = 12'h98F ;
assign kyber_zeta[18] = 12'h53B ;
assign kyber_zeta[19] = 12'h5C4 ;
assign kyber_zeta[20] = 12'hBE6 ;
assign kyber_zeta[21] = 12'h038 ;
assign kyber_zeta[22] = 12'h8C0 ;
assign kyber_zeta[23] = 12'h535 ;
assign kyber_zeta[24] = 12'h592 ;
assign kyber_zeta[25] = 12'h82E ;
assign kyber_zeta[26] = 12'h217 ;
assign kyber_zeta[27] = 12'hB42 ;
assign kyber_zeta[28] = 12'h959 ;
assign kyber_zeta[29] = 12'hB3F ;
assign kyber_zeta[30] = 12'h7B6 ;
assign kyber_zeta[31] = 12'h335 ;
assign kyber_zeta[32] = 12'h121 ;
assign kyber_zeta[33] = 12'h14B ;
assign kyber_zeta[34] = 12'hCB5 ;
assign kyber_zeta[35] = 12'h6DC ;
assign kyber_zeta[36] = 12'h4AD ;
assign kyber_zeta[37] = 12'h900 ;
assign kyber_zeta[38] = 12'h8E5 ;
assign kyber_zeta[39] = 12'h807 ;
assign kyber_zeta[40] = 12'h28A ;
assign kyber_zeta[41] = 12'h7B9 ;
assign kyber_zeta[42] = 12'h9D1 ;
assign kyber_zeta[43] = 12'h278 ;
assign kyber_zeta[44] = 12'hB31 ;
assign kyber_zeta[45] = 12'h021 ;
assign kyber_zeta[46] = 12'h528 ;
assign kyber_zeta[47] = 12'h77B ;
assign kyber_zeta[48] = 12'h90F ;
assign kyber_zeta[49] = 12'h59B ;
assign kyber_zeta[50] = 12'h327 ;
assign kyber_zeta[51] = 12'h1C4 ;
assign kyber_zeta[52] = 12'h59E ;
assign kyber_zeta[53] = 12'hB34 ;
assign kyber_zeta[54] = 12'h5FE ;
assign kyber_zeta[55] = 12'h962 ;
assign kyber_zeta[56] = 12'hA57 ;
assign kyber_zeta[57] = 12'hA39 ;
assign kyber_zeta[58] = 12'h5C9 ;
assign kyber_zeta[59] = 12'h288 ;
assign kyber_zeta[60] = 12'h9AA ;
assign kyber_zeta[61] = 12'hC26 ;
assign kyber_zeta[62] = 12'h4CB ;
assign kyber_zeta[63] = 12'h38E ;
assign kyber_zeta[64] = 12'h011 ;
assign kyber_zeta[65] = 12'hAC9 ;
assign kyber_zeta[66] = 12'h247 ;
assign kyber_zeta[67] = 12'hA59 ;
assign kyber_zeta[68] = 12'h665 ;
assign kyber_zeta[69] = 12'h2D3 ;
assign kyber_zeta[70] = 12'h8F0 ;
assign kyber_zeta[71] = 12'h44C ;
assign kyber_zeta[72] = 12'h581 ;
assign kyber_zeta[73] = 12'hA66 ;
assign kyber_zeta[74] = 12'hCD1 ;
assign kyber_zeta[75] = 12'h0E9 ;
assign kyber_zeta[76] = 12'h2F4 ;
assign kyber_zeta[77] = 12'h86C ;
assign kyber_zeta[78] = 12'hBC7 ;
assign kyber_zeta[79] = 12'hBEA ;
assign kyber_zeta[80] = 12'h6A7 ;
assign kyber_zeta[81] = 12'h673 ;
assign kyber_zeta[82] = 12'hAE5 ;
assign kyber_zeta[83] = 12'h6FD ;
assign kyber_zeta[84] = 12'h737 ;
assign kyber_zeta[85] = 12'h3B8 ;
assign kyber_zeta[86] = 12'h5B5 ;
assign kyber_zeta[87] = 12'hA7F ;
assign kyber_zeta[88] = 12'h3AB ;
assign kyber_zeta[89] = 12'h904 ;
assign kyber_zeta[90] = 12'h985 ;
assign kyber_zeta[91] = 12'h954 ;
assign kyber_zeta[92] = 12'h2DD ;
assign kyber_zeta[93] = 12'h921 ;
assign kyber_zeta[94] = 12'h10C ;
assign kyber_zeta[95] = 12'h281 ;
assign kyber_zeta[96] = 12'h630 ;
assign kyber_zeta[97] = 12'h8FA ;
assign kyber_zeta[98] = 12'h7F5 ;
assign kyber_zeta[99] = 12'hC94 ;
assign kyber_zeta[100] = 12'h177 ;
assign kyber_zeta[101] = 12'h9F5 ;
assign kyber_zeta[102] = 12'h82A ;
assign kyber_zeta[103] = 12'h66D ;
assign kyber_zeta[104] = 12'h427 ;
assign kyber_zeta[105] = 12'h13F ;
assign kyber_zeta[106] = 12'hAD5 ;
assign kyber_zeta[107] = 12'h2F5 ;
assign kyber_zeta[108] = 12'h833 ;
assign kyber_zeta[109] = 12'h231 ;
assign kyber_zeta[110] = 12'h9A2 ;
assign kyber_zeta[111] = 12'hA22 ;
assign kyber_zeta[112] = 12'hAF4 ;
assign kyber_zeta[113] = 12'h444 ;
assign kyber_zeta[114] = 12'h193 ;
assign kyber_zeta[115] = 12'h402 ;
assign kyber_zeta[116] = 12'h477 ;
assign kyber_zeta[117] = 12'h866 ;
assign kyber_zeta[118] = 12'hAD7 ;
assign kyber_zeta[119] = 12'h376 ;
assign kyber_zeta[120] = 12'h6BA ;
assign kyber_zeta[121] = 12'h4BC ;
assign kyber_zeta[122] = 12'h752 ;
assign kyber_zeta[123] = 12'h405 ;
assign kyber_zeta[124] = 12'h83E ;
assign kyber_zeta[125] = 12'hB77 ;
assign kyber_zeta[126] = 12'h375 ;
assign kyber_zeta[127] = 12'h86A ;
assign kyber_zeta[128] = 12'h011 ;
assign kyber_zeta[129] = 12'hCF0 ;
assign kyber_zeta[130] = 12'hAC9 ;
assign kyber_zeta[131] = 12'h238 ;
assign kyber_zeta[132] = 12'h247 ;
assign kyber_zeta[133] = 12'hABA ;
assign kyber_zeta[134] = 12'hA59 ;
assign kyber_zeta[135] = 12'h2A8 ;
assign kyber_zeta[136] = 12'h665 ;
assign kyber_zeta[137] = 12'h69C ;
assign kyber_zeta[138] = 12'h2D3 ;
assign kyber_zeta[139] = 12'hA2E ;
assign kyber_zeta[140] = 12'h8F0 ;
assign kyber_zeta[141] = 12'h411 ;
assign kyber_zeta[142] = 12'h44C ;
assign kyber_zeta[143] = 12'h8B5 ;
assign kyber_zeta[144] = 12'h581 ;
assign kyber_zeta[145] = 12'h780 ;
assign kyber_zeta[146] = 12'hA66 ;
assign kyber_zeta[147] = 12'h29B ;
assign kyber_zeta[148] = 12'hCD1 ;
assign kyber_zeta[149] = 12'h030 ;
assign kyber_zeta[150] = 12'h0E9 ;
assign kyber_zeta[151] = 12'hC18 ;
assign kyber_zeta[152] = 12'h2F4 ;
assign kyber_zeta[153] = 12'hA0D ;
assign kyber_zeta[154] = 12'h86C ;
assign kyber_zeta[155] = 12'h495 ;
assign kyber_zeta[156] = 12'hBC7 ;
assign kyber_zeta[157] = 12'h13A ;
assign kyber_zeta[158] = 12'hBEA ;
assign kyber_zeta[159] = 12'h117 ;
assign kyber_zeta[160] = 12'h6A7 ;
assign kyber_zeta[161] = 12'h65A ;
assign kyber_zeta[162] = 12'h673 ;
assign kyber_zeta[163] = 12'h68E ;
assign kyber_zeta[164] = 12'hAE5 ;
assign kyber_zeta[165] = 12'h21C ;
assign kyber_zeta[166] = 12'h6FD ;
assign kyber_zeta[167] = 12'h604 ;
assign kyber_zeta[168] = 12'h737 ;
assign kyber_zeta[169] = 12'h5CA ;
assign kyber_zeta[170] = 12'h3B8 ;
assign kyber_zeta[171] = 12'h949 ;
assign kyber_zeta[172] = 12'h5B5 ;
assign kyber_zeta[173] = 12'h74C ;
assign kyber_zeta[174] = 12'hA7F ;
assign kyber_zeta[175] = 12'h282 ;
assign kyber_zeta[176] = 12'h3AB ;
assign kyber_zeta[177] = 12'h956 ;
assign kyber_zeta[178] = 12'h904 ;
assign kyber_zeta[179] = 12'h3FD ;
assign kyber_zeta[180] = 12'h985 ;
assign kyber_zeta[181] = 12'h37C ;
assign kyber_zeta[182] = 12'h954 ;
assign kyber_zeta[183] = 12'h3AD ;
assign kyber_zeta[184] = 12'h2DD ;
assign kyber_zeta[185] = 12'hA24 ;
assign kyber_zeta[186] = 12'h921 ;
assign kyber_zeta[187] = 12'h3E0 ;
assign kyber_zeta[188] = 12'h10C ;
assign kyber_zeta[189] = 12'hBF5 ;
assign kyber_zeta[190] = 12'h281 ;
assign kyber_zeta[191] = 12'hA80 ;
assign kyber_zeta[192] = 12'h630 ;
assign kyber_zeta[193] = 12'h6D1 ;
assign kyber_zeta[194] = 12'h8FA ;
assign kyber_zeta[195] = 12'h407 ;
assign kyber_zeta[196] = 12'h7F5 ;
assign kyber_zeta[197] = 12'h50C ;
assign kyber_zeta[198] = 12'hC94 ;
assign kyber_zeta[199] = 12'h06D ;
assign kyber_zeta[200] = 12'h177 ;
assign kyber_zeta[201] = 12'hB8A ;
assign kyber_zeta[202] = 12'h9F5 ;
assign kyber_zeta[203] = 12'h30C ;
assign kyber_zeta[204] = 12'h82A ;
assign kyber_zeta[205] = 12'h4D7 ;
assign kyber_zeta[206] = 12'h66D ;
assign kyber_zeta[207] = 12'h694 ;
assign kyber_zeta[208] = 12'h427 ;
assign kyber_zeta[209] = 12'h8DA ;
assign kyber_zeta[210] = 12'h13F ;
assign kyber_zeta[211] = 12'hBC2 ;
assign kyber_zeta[212] = 12'hAD5 ;
assign kyber_zeta[213] = 12'h22C ;
assign kyber_zeta[214] = 12'h2F5 ;
assign kyber_zeta[215] = 12'hA0C ;
assign kyber_zeta[216] = 12'h833 ;
assign kyber_zeta[217] = 12'h4CE ;
assign kyber_zeta[218] = 12'h231 ;
assign kyber_zeta[219] = 12'hAD0 ;
assign kyber_zeta[220] = 12'h9A2 ;
assign kyber_zeta[221] = 12'h35F ;
assign kyber_zeta[222] = 12'hA22 ;
assign kyber_zeta[223] = 12'h2DF ;
assign kyber_zeta[224] = 12'hAF4 ;
assign kyber_zeta[225] = 12'h20D ;
assign kyber_zeta[226] = 12'h444 ;
assign kyber_zeta[227] = 12'h8BD ;
assign kyber_zeta[228] = 12'h193 ;
assign kyber_zeta[229] = 12'hB6E ;
assign kyber_zeta[230] = 12'h402 ;
assign kyber_zeta[231] = 12'h8FF ;
assign kyber_zeta[232] = 12'h477 ;
assign kyber_zeta[233] = 12'h88A ;
assign kyber_zeta[234] = 12'h866 ;
assign kyber_zeta[235] = 12'h49B ;
assign kyber_zeta[236] = 12'hAD7 ;
assign kyber_zeta[237] = 12'h22A ;
assign kyber_zeta[238] = 12'h376 ;
assign kyber_zeta[239] = 12'h98B ;
assign kyber_zeta[240] = 12'h6BA ;
assign kyber_zeta[241] = 12'h647 ;
assign kyber_zeta[242] = 12'h4BC ;
assign kyber_zeta[243] = 12'h845 ;
assign kyber_zeta[244] = 12'h752 ;
assign kyber_zeta[245] = 12'h5AF ;
assign kyber_zeta[246] = 12'h405 ;
assign kyber_zeta[247] = 12'h8FC ;
assign kyber_zeta[248] = 12'h83E ;
assign kyber_zeta[249] = 12'h4C3 ;
assign kyber_zeta[250] = 12'hB77 ;
assign kyber_zeta[251] = 12'h18A ;
assign kyber_zeta[252] = 12'h375 ;
assign kyber_zeta[253] = 12'h98C ;
assign kyber_zeta[254] = 12'h86A ;
assign kyber_zeta[255] = 12'h497 ;

//------------------------------------------------------------------------------------

assign kyber_zetainv[0] = 12'hD00 ;
assign kyber_zetainv[1] = 12'h640 ;
assign kyber_zetainv[2] = 12'h2ED ;
assign kyber_zetainv[3] = 12'h028 ;
assign kyber_zetainv[4] = 12'h2AF ;
assign kyber_zetainv[5] = 12'hA8B ;
assign kyber_zetainv[6] = 12'h598 ;
assign kyber_zetainv[7] = 12'h9B1 ;
assign kyber_zetainv[8] = 12'h8DB ;
assign kyber_zetainv[9] = 12'h582 ;
assign kyber_zetainv[10] = 12'hC40 ;
assign kyber_zetainv[11] = 12'h9E4 ;
assign kyber_zetainv[12] = 12'h21F ;
assign kyber_zetainv[13] = 12'h045 ;
assign kyber_zetainv[14] = 12'hAC8 ;
assign kyber_zetainv[15] = 12'h62F ;
assign kyber_zetainv[16] = 12'hBD9 ;
assign kyber_zetainv[17] = 12'h372 ;
assign kyber_zetainv[18] = 12'h7C6 ;
assign kyber_zetainv[19] = 12'h73D ;
assign kyber_zetainv[20] = 12'h11B ;
assign kyber_zetainv[21] = 12'hCC9 ;
assign kyber_zetainv[22] = 12'h441 ;
assign kyber_zetainv[23] = 12'h7CC ;
assign kyber_zetainv[24] = 12'h76F ;
assign kyber_zetainv[25] = 12'h4D3 ;
assign kyber_zetainv[26] = 12'hAEA ;
assign kyber_zetainv[27] = 12'h1BF ;
assign kyber_zetainv[28] = 12'h3A8 ;
assign kyber_zetainv[29] = 12'h1C2 ;
assign kyber_zetainv[30] = 12'h54B ;
assign kyber_zetainv[31] = 12'h9CC ;
assign kyber_zetainv[32] = 12'hBE0 ;
assign kyber_zetainv[33] = 12'hBB6 ;
assign kyber_zetainv[34] = 12'h04C ;
assign kyber_zetainv[35] = 12'h625 ;
assign kyber_zetainv[36] = 12'h854 ;
assign kyber_zetainv[37] = 12'h401 ;
assign kyber_zetainv[38] = 12'h41C ;
assign kyber_zetainv[39] = 12'h4FA ;
assign kyber_zetainv[40] = 12'hA77 ;
assign kyber_zetainv[41] = 12'h548 ;
assign kyber_zetainv[42] = 12'h330 ;
assign kyber_zetainv[43] = 12'hA89 ;
assign kyber_zetainv[44] = 12'h1D0 ;
assign kyber_zetainv[45] = 12'hCE0 ;
assign kyber_zetainv[46] = 12'h7D9 ;
assign kyber_zetainv[47] = 12'h586 ;
assign kyber_zetainv[48] = 12'h3F2 ;
assign kyber_zetainv[49] = 12'h766 ;
assign kyber_zetainv[50] = 12'h9DA ;
assign kyber_zetainv[51] = 12'hB3D ;
assign kyber_zetainv[52] = 12'h763 ;
assign kyber_zetainv[53] = 12'h1CD ;
assign kyber_zetainv[54] = 12'h703 ;
assign kyber_zetainv[55] = 12'h39F ;
assign kyber_zetainv[56] = 12'h2AA ;
assign kyber_zetainv[57] = 12'h2C8 ;
assign kyber_zetainv[58] = 12'h738 ;
assign kyber_zetainv[59] = 12'hA79 ;
assign kyber_zetainv[60] = 12'h357 ;
assign kyber_zetainv[61] = 12'h0DB ;
assign kyber_zetainv[62] = 12'h836 ;
assign kyber_zetainv[63] = 12'h973 ;
assign kyber_zetainv[64] = 12'hCF0 ;
assign kyber_zetainv[65] = 12'h238 ;
assign kyber_zetainv[66] = 12'hABA ;
assign kyber_zetainv[67] = 12'h2A8 ;
assign kyber_zetainv[68] = 12'h69C ;
assign kyber_zetainv[69] = 12'hA2E ;
assign kyber_zetainv[70] = 12'h411 ;
assign kyber_zetainv[71] = 12'h8B5 ;
assign kyber_zetainv[72] = 12'h780 ;
assign kyber_zetainv[73] = 12'h29B ;
assign kyber_zetainv[74] = 12'h030 ;
assign kyber_zetainv[75] = 12'hC18 ;
assign kyber_zetainv[76] = 12'hA0D ;
assign kyber_zetainv[77] = 12'h495 ;
assign kyber_zetainv[78] = 12'h13A ;
assign kyber_zetainv[79] = 12'h117 ;
assign kyber_zetainv[80] = 12'h65A ;
assign kyber_zetainv[81] = 12'h68E ;
assign kyber_zetainv[82] = 12'h21C ;
assign kyber_zetainv[83] = 12'h604 ;
assign kyber_zetainv[84] = 12'h5CA ;
assign kyber_zetainv[85] = 12'h949 ;
assign kyber_zetainv[86] = 12'h74C ;
assign kyber_zetainv[87] = 12'h282 ;
assign kyber_zetainv[88] = 12'h956 ;
assign kyber_zetainv[89] = 12'h3FD ;
assign kyber_zetainv[90] = 12'h37C ;
assign kyber_zetainv[91] = 12'h3AD ;
assign kyber_zetainv[92] = 12'hA24 ;
assign kyber_zetainv[93] = 12'h3E0 ;
assign kyber_zetainv[94] = 12'hBF5 ;
assign kyber_zetainv[95] = 12'hA80 ;
assign kyber_zetainv[96] = 12'h6D1 ;
assign kyber_zetainv[97] = 12'h407 ;
assign kyber_zetainv[98] = 12'h50C ;
assign kyber_zetainv[99] = 12'h06D ;
assign kyber_zetainv[100] = 12'hB8A ;
assign kyber_zetainv[101] = 12'h30C ;
assign kyber_zetainv[102] = 12'h4D7 ;
assign kyber_zetainv[103] = 12'h694 ;
assign kyber_zetainv[104] = 12'h8DA ;
assign kyber_zetainv[105] = 12'hBC2 ;
assign kyber_zetainv[106] = 12'h22C ;
assign kyber_zetainv[107] = 12'hA0C ;
assign kyber_zetainv[108] = 12'h4CE ;
assign kyber_zetainv[109] = 12'hAD0 ;
assign kyber_zetainv[110] = 12'h35F ;
assign kyber_zetainv[111] = 12'h2DF ;
assign kyber_zetainv[112] = 12'h20D ;
assign kyber_zetainv[113] = 12'h8BD ;
assign kyber_zetainv[114] = 12'hB6E ;
assign kyber_zetainv[115] = 12'h8FF ;
assign kyber_zetainv[116] = 12'h88A ;
assign kyber_zetainv[117] = 12'h49B ;
assign kyber_zetainv[118] = 12'h22A ;
assign kyber_zetainv[119] = 12'h98B ;
assign kyber_zetainv[120] = 12'h647 ;
assign kyber_zetainv[121] = 12'h845 ;
assign kyber_zetainv[122] = 12'h5AF ;
assign kyber_zetainv[123] = 12'h8FC ;
assign kyber_zetainv[124] = 12'h4C3 ;
assign kyber_zetainv[125] = 12'h18A ;
assign kyber_zetainv[126] = 12'h98C ;
assign kyber_zetainv[127] = 12'h497 ;
assign kyber_zetainv[128] = 12'hCF0 ;
assign kyber_zetainv[129] = 12'h011 ;
assign kyber_zetainv[130] = 12'h238 ;
assign kyber_zetainv[131] = 12'hAC9 ;
assign kyber_zetainv[132] = 12'hABA ;
assign kyber_zetainv[133] = 12'h247 ;
assign kyber_zetainv[134] = 12'h2A8 ;
assign kyber_zetainv[135] = 12'hA59 ;
assign kyber_zetainv[136] = 12'h69C ;
assign kyber_zetainv[137] = 12'h665 ;
assign kyber_zetainv[138] = 12'hA2E ;
assign kyber_zetainv[139] = 12'h2D3 ;
assign kyber_zetainv[140] = 12'h411 ;
assign kyber_zetainv[141] = 12'h8F0 ;
assign kyber_zetainv[142] = 12'h8B5 ;
assign kyber_zetainv[143] = 12'h44C ;
assign kyber_zetainv[144] = 12'h780 ;
assign kyber_zetainv[145] = 12'h581 ;
assign kyber_zetainv[146] = 12'h29B ;
assign kyber_zetainv[147] = 12'hA66 ;
assign kyber_zetainv[148] = 12'h030 ;
assign kyber_zetainv[149] = 12'hCD1 ;
assign kyber_zetainv[150] = 12'hC18 ;
assign kyber_zetainv[151] = 12'h0E9 ;
assign kyber_zetainv[152] = 12'hA0D ;
assign kyber_zetainv[153] = 12'h2F4 ;
assign kyber_zetainv[154] = 12'h495 ;
assign kyber_zetainv[155] = 12'h86C ;
assign kyber_zetainv[156] = 12'h13A ;
assign kyber_zetainv[157] = 12'hBC7 ;
assign kyber_zetainv[158] = 12'h117 ;
assign kyber_zetainv[159] = 12'hBEA ;
assign kyber_zetainv[160] = 12'h65A ;
assign kyber_zetainv[161] = 12'h6A7 ;
assign kyber_zetainv[162] = 12'h68E ;
assign kyber_zetainv[163] = 12'h673 ;
assign kyber_zetainv[164] = 12'h21C ;
assign kyber_zetainv[165] = 12'hAE5 ;
assign kyber_zetainv[166] = 12'h604 ;
assign kyber_zetainv[167] = 12'h6FD ;
assign kyber_zetainv[168] = 12'h5CA ;
assign kyber_zetainv[169] = 12'h737 ;
assign kyber_zetainv[170] = 12'h949 ;
assign kyber_zetainv[171] = 12'h3B8 ;
assign kyber_zetainv[172] = 12'h74C ;
assign kyber_zetainv[173] = 12'h5B5 ;
assign kyber_zetainv[174] = 12'h282 ;
assign kyber_zetainv[175] = 12'hA7F ;
assign kyber_zetainv[176] = 12'h956 ;
assign kyber_zetainv[177] = 12'h3AB ;
assign kyber_zetainv[178] = 12'h3FD ;
assign kyber_zetainv[179] = 12'h904 ;
assign kyber_zetainv[180] = 12'h37C ;
assign kyber_zetainv[181] = 12'h985 ;
assign kyber_zetainv[182] = 12'h3AD ;
assign kyber_zetainv[183] = 12'h954 ;
assign kyber_zetainv[184] = 12'hA24 ;
assign kyber_zetainv[185] = 12'h2DD ;
assign kyber_zetainv[186] = 12'h3E0 ;
assign kyber_zetainv[187] = 12'h921 ;
assign kyber_zetainv[188] = 12'hBF5 ;
assign kyber_zetainv[189] = 12'h10C ;
assign kyber_zetainv[190] = 12'hA80 ;
assign kyber_zetainv[191] = 12'h281 ;
assign kyber_zetainv[192] = 12'h6D1 ;
assign kyber_zetainv[193] = 12'h630 ;
assign kyber_zetainv[194] = 12'h407 ;
assign kyber_zetainv[195] = 12'h8FA ;
assign kyber_zetainv[196] = 12'h50C ;
assign kyber_zetainv[197] = 12'h7F5 ;
assign kyber_zetainv[198] = 12'h06D ;
assign kyber_zetainv[199] = 12'hC94 ;
assign kyber_zetainv[200] = 12'hB8A ;
assign kyber_zetainv[201] = 12'h177 ;
assign kyber_zetainv[202] = 12'h30C ;
assign kyber_zetainv[203] = 12'h9F5 ;
assign kyber_zetainv[204] = 12'h4D7 ;
assign kyber_zetainv[205] = 12'h82A ;
assign kyber_zetainv[206] = 12'h694 ;
assign kyber_zetainv[207] = 12'h66D ;
assign kyber_zetainv[208] = 12'h8DA ;
assign kyber_zetainv[209] = 12'h427 ;
assign kyber_zetainv[210] = 12'hBC2 ;
assign kyber_zetainv[211] = 12'h13F ;
assign kyber_zetainv[212] = 12'h22C ;
assign kyber_zetainv[213] = 12'hAD5 ;
assign kyber_zetainv[214] = 12'hA0C ;
assign kyber_zetainv[215] = 12'h2F5 ;
assign kyber_zetainv[216] = 12'h4CE ;
assign kyber_zetainv[217] = 12'h833 ;
assign kyber_zetainv[218] = 12'hAD0 ;
assign kyber_zetainv[219] = 12'h231 ;
assign kyber_zetainv[220] = 12'h35F ;
assign kyber_zetainv[221] = 12'h9A2 ;
assign kyber_zetainv[222] = 12'h2DF ;
assign kyber_zetainv[223] = 12'hA22 ;
assign kyber_zetainv[224] = 12'h20D ;
assign kyber_zetainv[225] = 12'hAF4 ;
assign kyber_zetainv[226] = 12'h8BD ;
assign kyber_zetainv[227] = 12'h444 ;
assign kyber_zetainv[228] = 12'hB6E ;
assign kyber_zetainv[229] = 12'h193 ;
assign kyber_zetainv[230] = 12'h8FF ;
assign kyber_zetainv[231] = 12'h402 ;
assign kyber_zetainv[232] = 12'h88A ;
assign kyber_zetainv[233] = 12'h477 ;
assign kyber_zetainv[234] = 12'h49B ;
assign kyber_zetainv[235] = 12'h866 ;
assign kyber_zetainv[236] = 12'h22A ;
assign kyber_zetainv[237] = 12'hAD7 ;
assign kyber_zetainv[238] = 12'h98B ;
assign kyber_zetainv[239] = 12'h376 ;
assign kyber_zetainv[240] = 12'h647 ;
assign kyber_zetainv[241] = 12'h6BA ;
assign kyber_zetainv[242] = 12'h845 ;
assign kyber_zetainv[243] = 12'h4BC ;
assign kyber_zetainv[244] = 12'h5AF ;
assign kyber_zetainv[245] = 12'h752 ;
assign kyber_zetainv[246] = 12'h8FC ;
assign kyber_zetainv[247] = 12'h405 ;
assign kyber_zetainv[248] = 12'h4C3 ;
assign kyber_zetainv[249] = 12'h83E ;
assign kyber_zetainv[250] = 12'h18A ;
assign kyber_zetainv[251] = 12'hB77 ;
assign kyber_zetainv[252] = 12'h98C ;
assign kyber_zetainv[253] = 12'h375 ;
assign kyber_zetainv[254] = 12'h497 ;
assign kyber_zetainv[255] = 12'h86A ;

// assign ntt_twiddle_mem[0]  = 'h000001;
assign ntt_twiddle_mem[0]  = {zeta[3],  zeta[2],  zeta[1]};
assign ntt_twiddle_mem[1]  = {zeta[9],  zeta[8],  zeta[4]};
assign ntt_twiddle_mem[2]  = {zeta[11], zeta[10], zeta[5]};
assign ntt_twiddle_mem[3]  = {zeta[13], zeta[12], zeta[6]};
assign ntt_twiddle_mem[4]  = {zeta[15], zeta[14], zeta[7]};
assign ntt_twiddle_mem[5]  = {zeta[33], zeta[32], zeta[16]};
assign ntt_twiddle_mem[6]  = {zeta[35], zeta[34], zeta[17]};
assign ntt_twiddle_mem[7]  = {zeta[37], zeta[36], zeta[18]};
assign ntt_twiddle_mem[8]  = {zeta[39], zeta[38], zeta[19]};
assign ntt_twiddle_mem[9]  = {zeta[41], zeta[40], zeta[20]};
assign ntt_twiddle_mem[10] = {zeta[43], zeta[42], zeta[21]};
assign ntt_twiddle_mem[11] = {zeta[45], zeta[44], zeta[22]};
assign ntt_twiddle_mem[12] = {zeta[47], zeta[46], zeta[23]};
assign ntt_twiddle_mem[13] = {zeta[49], zeta[48], zeta[24]};
assign ntt_twiddle_mem[14] = {zeta[51], zeta[50], zeta[25]};
assign ntt_twiddle_mem[15] = {zeta[53], zeta[52], zeta[26]};
assign ntt_twiddle_mem[16] = {zeta[55], zeta[54], zeta[27]};
assign ntt_twiddle_mem[17] = {zeta[57], zeta[56], zeta[28]};
assign ntt_twiddle_mem[18] = {zeta[59], zeta[58], zeta[29]};
assign ntt_twiddle_mem[19] = {zeta[61], zeta[60], zeta[30]};
assign ntt_twiddle_mem[20] = {zeta[63], zeta[62], zeta[31]};
assign ntt_twiddle_mem[21] = {zeta[129], zeta[128], zeta[64]};
assign ntt_twiddle_mem[22] = {zeta[131], zeta[130], zeta[65]};
assign ntt_twiddle_mem[23] = {zeta[133], zeta[132], zeta[66]};
assign ntt_twiddle_mem[24] = {zeta[135], zeta[134], zeta[67]};
assign ntt_twiddle_mem[25] = {zeta[137], zeta[136], zeta[68]};
assign ntt_twiddle_mem[26] = {zeta[139], zeta[138], zeta[69]};
assign ntt_twiddle_mem[27] = {zeta[141], zeta[140], zeta[70]};
assign ntt_twiddle_mem[28] = {zeta[143], zeta[142], zeta[71]};
assign ntt_twiddle_mem[29] = {zeta[145], zeta[144], zeta[72]};
assign ntt_twiddle_mem[30] = {zeta[147], zeta[146], zeta[73]};
assign ntt_twiddle_mem[31] = {zeta[149], zeta[148], zeta[74]};
assign ntt_twiddle_mem[32] = {zeta[151], zeta[150], zeta[75]};
assign ntt_twiddle_mem[33] = {zeta[153], zeta[152], zeta[76]};
assign ntt_twiddle_mem[34] = {zeta[155], zeta[154], zeta[77]};
assign ntt_twiddle_mem[35] = {zeta[157], zeta[156], zeta[78]};
assign ntt_twiddle_mem[36] = {zeta[159], zeta[158], zeta[79]};
assign ntt_twiddle_mem[37] = {zeta[161], zeta[160], zeta[80]};
assign ntt_twiddle_mem[38] = {zeta[163], zeta[162], zeta[81]};
assign ntt_twiddle_mem[39] = {zeta[165], zeta[164], zeta[82]};
assign ntt_twiddle_mem[40] = {zeta[167], zeta[166], zeta[83]};
assign ntt_twiddle_mem[41] = {zeta[169], zeta[168], zeta[84]};
assign ntt_twiddle_mem[42] = {zeta[171], zeta[170], zeta[85]};
assign ntt_twiddle_mem[43] = {zeta[173], zeta[172], zeta[86]};
assign ntt_twiddle_mem[44] = {zeta[175], zeta[174], zeta[87]};
assign ntt_twiddle_mem[45] = {zeta[177], zeta[176], zeta[88]};
assign ntt_twiddle_mem[46] = {zeta[179], zeta[178], zeta[89]};
assign ntt_twiddle_mem[47] = {zeta[181], zeta[180], zeta[90]};
assign ntt_twiddle_mem[48] = {zeta[183], zeta[182], zeta[91]};
assign ntt_twiddle_mem[49] = {zeta[185], zeta[184], zeta[92]};
assign ntt_twiddle_mem[50] = {zeta[187], zeta[186], zeta[93]};
assign ntt_twiddle_mem[51] = {zeta[189], zeta[188], zeta[94]};
assign ntt_twiddle_mem[52] = {zeta[191], zeta[190], zeta[95]};
assign ntt_twiddle_mem[53] = {zeta[193], zeta[192], zeta[96]};
assign ntt_twiddle_mem[54] = {zeta[195], zeta[194], zeta[97]};
assign ntt_twiddle_mem[55] = {zeta[197], zeta[196], zeta[98]};
assign ntt_twiddle_mem[56] = {zeta[199], zeta[198], zeta[99]};
assign ntt_twiddle_mem[57] = {zeta[201], zeta[200], zeta[100]};
assign ntt_twiddle_mem[58] = {zeta[203], zeta[202], zeta[101]};
assign ntt_twiddle_mem[59] = {zeta[205], zeta[204], zeta[102]};
assign ntt_twiddle_mem[60] = {zeta[207], zeta[206], zeta[103]};
assign ntt_twiddle_mem[61] = {zeta[209], zeta[208], zeta[104]};
assign ntt_twiddle_mem[62] = {zeta[211], zeta[210], zeta[105]};
assign ntt_twiddle_mem[63] = {zeta[213], zeta[212], zeta[106]};
assign ntt_twiddle_mem[64] = {zeta[215], zeta[214], zeta[107]};
assign ntt_twiddle_mem[65] = {zeta[217], zeta[216], zeta[108]};
assign ntt_twiddle_mem[66] = {zeta[219], zeta[218], zeta[109]};
assign ntt_twiddle_mem[67] = {zeta[221], zeta[220], zeta[110]};
assign ntt_twiddle_mem[68] = {zeta[223], zeta[222], zeta[111]};
assign ntt_twiddle_mem[69] = {zeta[225], zeta[224], zeta[112]};
assign ntt_twiddle_mem[70] = {zeta[227], zeta[226], zeta[113]};
assign ntt_twiddle_mem[71] = {zeta[229], zeta[228], zeta[114]};
assign ntt_twiddle_mem[72] = {zeta[231], zeta[230], zeta[115]};
assign ntt_twiddle_mem[73] = {zeta[233], zeta[232], zeta[116]};
assign ntt_twiddle_mem[74] = {zeta[235], zeta[234], zeta[117]};
assign ntt_twiddle_mem[75] = {zeta[237], zeta[236], zeta[118]};
assign ntt_twiddle_mem[76] = {zeta[239], zeta[238], zeta[119]};
assign ntt_twiddle_mem[77] = {zeta[241], zeta[240], zeta[120]};
assign ntt_twiddle_mem[78] = {zeta[243], zeta[242], zeta[121]};
assign ntt_twiddle_mem[79] = {zeta[245], zeta[244], zeta[122]};
assign ntt_twiddle_mem[80] = {zeta[247], zeta[246], zeta[123]};
assign ntt_twiddle_mem[81] = {zeta[249], zeta[248], zeta[124]};
assign ntt_twiddle_mem[82] = {zeta[251], zeta[250], zeta[125]};
assign ntt_twiddle_mem[83] = {zeta[253], zeta[252], zeta[126]};
assign ntt_twiddle_mem[84] = {zeta[255], zeta[254], zeta[127]};
//--------------------------------------------------------

assign intt_twiddle_mem[0]  = {zetainv[127], zetainv[254], zetainv[255]};
assign intt_twiddle_mem[1]  = {zetainv[126], zetainv[252], zetainv[253]};
assign intt_twiddle_mem[2]  = {zetainv[125], zetainv[250], zetainv[251]};
assign intt_twiddle_mem[3]  = {zetainv[124], zetainv[248], zetainv[249]};
assign intt_twiddle_mem[4]  = {zetainv[123], zetainv[246], zetainv[247]};
assign intt_twiddle_mem[5]  = {zetainv[122], zetainv[244], zetainv[245]};
assign intt_twiddle_mem[6]  = {zetainv[121], zetainv[242], zetainv[243]};
assign intt_twiddle_mem[7]  = {zetainv[120], zetainv[240], zetainv[241]};
assign intt_twiddle_mem[8]  = {zetainv[119], zetainv[238], zetainv[239]};
assign intt_twiddle_mem[9]  = {zetainv[118], zetainv[236], zetainv[237]};
assign intt_twiddle_mem[10] = {zetainv[117], zetainv[234], zetainv[235]};
assign intt_twiddle_mem[11] = {zetainv[116], zetainv[232], zetainv[233]};
assign intt_twiddle_mem[12] = {zetainv[115], zetainv[230], zetainv[231]};
assign intt_twiddle_mem[13] = {zetainv[114], zetainv[228], zetainv[229]};
assign intt_twiddle_mem[14] = {zetainv[113], zetainv[226], zetainv[227]};
assign intt_twiddle_mem[15] = {zetainv[112], zetainv[224], zetainv[225]};
assign intt_twiddle_mem[16] = {zetainv[111], zetainv[222], zetainv[223]};
assign intt_twiddle_mem[17] = {zetainv[110], zetainv[220], zetainv[221]};
assign intt_twiddle_mem[18] = {zetainv[109], zetainv[218], zetainv[219]};
assign intt_twiddle_mem[19] = {zetainv[108], zetainv[216], zetainv[217]};
assign intt_twiddle_mem[20] = {zetainv[107], zetainv[214], zetainv[215]};
assign intt_twiddle_mem[21] = {zetainv[106], zetainv[212], zetainv[213]};
assign intt_twiddle_mem[22] = {zetainv[105], zetainv[210], zetainv[211]};
assign intt_twiddle_mem[23] = {zetainv[104], zetainv[208], zetainv[209]};
assign intt_twiddle_mem[24] = {zetainv[103], zetainv[206], zetainv[207]};
assign intt_twiddle_mem[25] = {zetainv[102], zetainv[204], zetainv[205]};
assign intt_twiddle_mem[26] = {zetainv[101], zetainv[202], zetainv[203]};
assign intt_twiddle_mem[27] = {zetainv[100], zetainv[200], zetainv[201]};
assign intt_twiddle_mem[28] = {zetainv[99], zetainv[198], zetainv[199]};
assign intt_twiddle_mem[29] = {zetainv[98], zetainv[196], zetainv[197]};
assign intt_twiddle_mem[30] = {zetainv[97], zetainv[194], zetainv[195]};
assign intt_twiddle_mem[31] = {zetainv[96], zetainv[192], zetainv[193]};
assign intt_twiddle_mem[32] = {zetainv[95], zetainv[190], zetainv[191]};
assign intt_twiddle_mem[33] = {zetainv[94], zetainv[188], zetainv[189]};
assign intt_twiddle_mem[34] = {zetainv[93], zetainv[186], zetainv[187]};
assign intt_twiddle_mem[35] = {zetainv[92], zetainv[184], zetainv[185]};
assign intt_twiddle_mem[36] = {zetainv[91], zetainv[182], zetainv[183]};
assign intt_twiddle_mem[37] = {zetainv[90], zetainv[180], zetainv[181]};
assign intt_twiddle_mem[38] = {zetainv[89], zetainv[178], zetainv[179]};
assign intt_twiddle_mem[39] = {zetainv[88], zetainv[176], zetainv[177]};
assign intt_twiddle_mem[40] = {zetainv[87], zetainv[174], zetainv[175]};
assign intt_twiddle_mem[41] = {zetainv[86], zetainv[172], zetainv[173]};
assign intt_twiddle_mem[42] = {zetainv[85], zetainv[170], zetainv[171]};
assign intt_twiddle_mem[43] = {zetainv[84], zetainv[168], zetainv[169]};
assign intt_twiddle_mem[44] = {zetainv[83], zetainv[166], zetainv[167]};
assign intt_twiddle_mem[45] = {zetainv[82], zetainv[164], zetainv[165]};
assign intt_twiddle_mem[46] = {zetainv[81], zetainv[162], zetainv[163]};
assign intt_twiddle_mem[47] = {zetainv[80], zetainv[160], zetainv[161]};
assign intt_twiddle_mem[48] = {zetainv[79], zetainv[158], zetainv[159]};
assign intt_twiddle_mem[49] = {zetainv[78], zetainv[156], zetainv[157]};
assign intt_twiddle_mem[50] = {zetainv[77], zetainv[154], zetainv[155]};
assign intt_twiddle_mem[51] = {zetainv[76], zetainv[152], zetainv[153]};
assign intt_twiddle_mem[52] = {zetainv[75], zetainv[150], zetainv[151]};
assign intt_twiddle_mem[53] = {zetainv[74], zetainv[148], zetainv[149]};
assign intt_twiddle_mem[54] = {zetainv[73], zetainv[146], zetainv[147]};
assign intt_twiddle_mem[55] = {zetainv[72], zetainv[144], zetainv[145]};
assign intt_twiddle_mem[56] = {zetainv[71], zetainv[142], zetainv[143]};
assign intt_twiddle_mem[57] = {zetainv[70], zetainv[140], zetainv[141]};
assign intt_twiddle_mem[58] = {zetainv[69], zetainv[138], zetainv[139]};
assign intt_twiddle_mem[59] = {zetainv[68], zetainv[136], zetainv[137]};
assign intt_twiddle_mem[60] = {zetainv[67], zetainv[134], zetainv[135]};
assign intt_twiddle_mem[61] = {zetainv[66], zetainv[132], zetainv[133]};
assign intt_twiddle_mem[62] = {zetainv[65], zetainv[130], zetainv[131]};
assign intt_twiddle_mem[63] = {zetainv[64], zetainv[128], zetainv[129]};
assign intt_twiddle_mem[64] = {zetainv[31], zetainv[62], zetainv[63]};
assign intt_twiddle_mem[65] = {zetainv[30], zetainv[60], zetainv[61]};
assign intt_twiddle_mem[66] = {zetainv[29], zetainv[58], zetainv[59]}; 
assign intt_twiddle_mem[67] = {zetainv[28], zetainv[56], zetainv[57]};
assign intt_twiddle_mem[68] = {zetainv[27], zetainv[54], zetainv[55]};
assign intt_twiddle_mem[69] = {zetainv[26], zetainv[52], zetainv[53]};
assign intt_twiddle_mem[70] = {zetainv[25], zetainv[50], zetainv[51]};
assign intt_twiddle_mem[71] = {zetainv[24], zetainv[48], zetainv[49]};
assign intt_twiddle_mem[72] = {zetainv[23], zetainv[46], zetainv[47]};
assign intt_twiddle_mem[73] = {zetainv[22], zetainv[44], zetainv[45]};
assign intt_twiddle_mem[74] = {zetainv[21], zetainv[42], zetainv[43]};
assign intt_twiddle_mem[75] = {zetainv[20], zetainv[40], zetainv[41]};
assign intt_twiddle_mem[76] = {zetainv[19], zetainv[38], zetainv[39]};
assign intt_twiddle_mem[77] = {zetainv[18], zetainv[36], zetainv[37]};
assign intt_twiddle_mem[78] = {zetainv[17], zetainv[34], zetainv[35]};
assign intt_twiddle_mem[79] = {zetainv[16], zetainv[32], zetainv[33]};
assign intt_twiddle_mem[80] = {zetainv[7], zetainv[14], zetainv[15]};
assign intt_twiddle_mem[81] = {zetainv[6], zetainv[12], zetainv[13]};
assign intt_twiddle_mem[82] = {zetainv[5], zetainv[10], zetainv[11]};
assign intt_twiddle_mem[83] = {zetainv[4], zetainv[8], zetainv[9]};
assign intt_twiddle_mem[84] = {zetainv[1], zetainv[2], zetainv[3]};

//--------------------------------------------------------

assign kyber_ntt_twiddle_mem[0]  = {kyber_zeta[3],  kyber_zeta[2],  kyber_zeta[1]};
assign kyber_ntt_twiddle_mem[1]  = {kyber_zeta[9],  kyber_zeta[8],  kyber_zeta[4]};
assign kyber_ntt_twiddle_mem[2]  = {kyber_zeta[11], kyber_zeta[10], kyber_zeta[5]};
assign kyber_ntt_twiddle_mem[3]  = {kyber_zeta[13], kyber_zeta[12], kyber_zeta[6]};
assign kyber_ntt_twiddle_mem[4]  = {kyber_zeta[15], kyber_zeta[14], kyber_zeta[7]};
assign kyber_ntt_twiddle_mem[5]  = {kyber_zeta[33], kyber_zeta[32], kyber_zeta[16]};
assign kyber_ntt_twiddle_mem[6]  = {kyber_zeta[35], kyber_zeta[34], kyber_zeta[17]};
assign kyber_ntt_twiddle_mem[7]  = {kyber_zeta[37], kyber_zeta[36], kyber_zeta[18]};
assign kyber_ntt_twiddle_mem[8]  = {kyber_zeta[39], kyber_zeta[38], kyber_zeta[19]};
assign kyber_ntt_twiddle_mem[9]  = {kyber_zeta[41], kyber_zeta[40], kyber_zeta[20]};
assign kyber_ntt_twiddle_mem[10] = {kyber_zeta[43], kyber_zeta[42], kyber_zeta[21]};
assign kyber_ntt_twiddle_mem[11] = {kyber_zeta[45], kyber_zeta[44], kyber_zeta[22]};
assign kyber_ntt_twiddle_mem[12] = {kyber_zeta[47], kyber_zeta[46], kyber_zeta[23]};
assign kyber_ntt_twiddle_mem[13] = {kyber_zeta[49], kyber_zeta[48], kyber_zeta[24]};
assign kyber_ntt_twiddle_mem[14] = {kyber_zeta[51], kyber_zeta[50], kyber_zeta[25]};
assign kyber_ntt_twiddle_mem[15] = {kyber_zeta[53], kyber_zeta[52], kyber_zeta[26]};
assign kyber_ntt_twiddle_mem[16] = {kyber_zeta[55], kyber_zeta[54], kyber_zeta[27]};
assign kyber_ntt_twiddle_mem[17] = {kyber_zeta[57], kyber_zeta[56], kyber_zeta[28]};
assign kyber_ntt_twiddle_mem[18] = {kyber_zeta[59], kyber_zeta[58], kyber_zeta[29]};
assign kyber_ntt_twiddle_mem[19] = {kyber_zeta[61], kyber_zeta[60], kyber_zeta[30]};
assign kyber_ntt_twiddle_mem[20] = {kyber_zeta[63], kyber_zeta[62], kyber_zeta[31]};
assign kyber_ntt_twiddle_mem[21] = {kyber_zeta[129], kyber_zeta[128], kyber_zeta[64]};
assign kyber_ntt_twiddle_mem[22] = {kyber_zeta[131], kyber_zeta[130], kyber_zeta[65]};
assign kyber_ntt_twiddle_mem[23] = {kyber_zeta[133], kyber_zeta[132], kyber_zeta[66]};
assign kyber_ntt_twiddle_mem[24] = {kyber_zeta[135], kyber_zeta[134], kyber_zeta[67]};
assign kyber_ntt_twiddle_mem[25] = {kyber_zeta[137], kyber_zeta[136], kyber_zeta[68]};
assign kyber_ntt_twiddle_mem[26] = {kyber_zeta[139], kyber_zeta[138], kyber_zeta[69]};
assign kyber_ntt_twiddle_mem[27] = {kyber_zeta[141], kyber_zeta[140], kyber_zeta[70]};
assign kyber_ntt_twiddle_mem[28] = {kyber_zeta[143], kyber_zeta[142], kyber_zeta[71]};
assign kyber_ntt_twiddle_mem[29] = {kyber_zeta[145], kyber_zeta[144], kyber_zeta[72]};
assign kyber_ntt_twiddle_mem[30] = {kyber_zeta[147], kyber_zeta[146], kyber_zeta[73]};
assign kyber_ntt_twiddle_mem[31] = {kyber_zeta[149], kyber_zeta[148], kyber_zeta[74]};
assign kyber_ntt_twiddle_mem[32] = {kyber_zeta[151], kyber_zeta[150], kyber_zeta[75]};
assign kyber_ntt_twiddle_mem[33] = {kyber_zeta[153], kyber_zeta[152], kyber_zeta[76]};
assign kyber_ntt_twiddle_mem[34] = {kyber_zeta[155], kyber_zeta[154], kyber_zeta[77]};
assign kyber_ntt_twiddle_mem[35] = {kyber_zeta[157], kyber_zeta[156], kyber_zeta[78]};
assign kyber_ntt_twiddle_mem[36] = {kyber_zeta[159], kyber_zeta[158], kyber_zeta[79]};
assign kyber_ntt_twiddle_mem[37] = {kyber_zeta[161], kyber_zeta[160], kyber_zeta[80]};
assign kyber_ntt_twiddle_mem[38] = {kyber_zeta[163], kyber_zeta[162], kyber_zeta[81]};
assign kyber_ntt_twiddle_mem[39] = {kyber_zeta[165], kyber_zeta[164], kyber_zeta[82]};
assign kyber_ntt_twiddle_mem[40] = {kyber_zeta[167], kyber_zeta[166], kyber_zeta[83]};
assign kyber_ntt_twiddle_mem[41] = {kyber_zeta[169], kyber_zeta[168], kyber_zeta[84]};
assign kyber_ntt_twiddle_mem[42] = {kyber_zeta[171], kyber_zeta[170], kyber_zeta[85]};
assign kyber_ntt_twiddle_mem[43] = {kyber_zeta[173], kyber_zeta[172], kyber_zeta[86]};
assign kyber_ntt_twiddle_mem[44] = {kyber_zeta[175], kyber_zeta[174], kyber_zeta[87]};
assign kyber_ntt_twiddle_mem[45] = {kyber_zeta[177], kyber_zeta[176], kyber_zeta[88]};
assign kyber_ntt_twiddle_mem[46] = {kyber_zeta[179], kyber_zeta[178], kyber_zeta[89]};
assign kyber_ntt_twiddle_mem[47] = {kyber_zeta[181], kyber_zeta[180], kyber_zeta[90]};
assign kyber_ntt_twiddle_mem[48] = {kyber_zeta[183], kyber_zeta[182], kyber_zeta[91]};
assign kyber_ntt_twiddle_mem[49] = {kyber_zeta[185], kyber_zeta[184], kyber_zeta[92]};
assign kyber_ntt_twiddle_mem[50] = {kyber_zeta[187], kyber_zeta[186], kyber_zeta[93]};
assign kyber_ntt_twiddle_mem[51] = {kyber_zeta[189], kyber_zeta[188], kyber_zeta[94]};
assign kyber_ntt_twiddle_mem[52] = {kyber_zeta[191], kyber_zeta[190], kyber_zeta[95]};
assign kyber_ntt_twiddle_mem[53] = {kyber_zeta[193], kyber_zeta[192], kyber_zeta[96]};
assign kyber_ntt_twiddle_mem[54] = {kyber_zeta[195], kyber_zeta[194], kyber_zeta[97]};
assign kyber_ntt_twiddle_mem[55] = {kyber_zeta[197], kyber_zeta[196], kyber_zeta[98]};
assign kyber_ntt_twiddle_mem[56] = {kyber_zeta[199], kyber_zeta[198], kyber_zeta[99]};
assign kyber_ntt_twiddle_mem[57] = {kyber_zeta[201], kyber_zeta[200], kyber_zeta[100]};
assign kyber_ntt_twiddle_mem[58] = {kyber_zeta[203], kyber_zeta[202], kyber_zeta[101]};
assign kyber_ntt_twiddle_mem[59] = {kyber_zeta[205], kyber_zeta[204], kyber_zeta[102]};
assign kyber_ntt_twiddle_mem[60] = {kyber_zeta[207], kyber_zeta[206], kyber_zeta[103]};
assign kyber_ntt_twiddle_mem[61] = {kyber_zeta[209], kyber_zeta[208], kyber_zeta[104]};
assign kyber_ntt_twiddle_mem[62] = {kyber_zeta[211], kyber_zeta[210], kyber_zeta[105]};
assign kyber_ntt_twiddle_mem[63] = {kyber_zeta[213], kyber_zeta[212], kyber_zeta[106]};
assign kyber_ntt_twiddle_mem[64] = {kyber_zeta[215], kyber_zeta[214], kyber_zeta[107]};
assign kyber_ntt_twiddle_mem[65] = {kyber_zeta[217], kyber_zeta[216], kyber_zeta[108]};
assign kyber_ntt_twiddle_mem[66] = {kyber_zeta[219], kyber_zeta[218], kyber_zeta[109]};
assign kyber_ntt_twiddle_mem[67] = {kyber_zeta[221], kyber_zeta[220], kyber_zeta[110]};
assign kyber_ntt_twiddle_mem[68] = {kyber_zeta[223], kyber_zeta[222], kyber_zeta[111]};
assign kyber_ntt_twiddle_mem[69] = {kyber_zeta[225], kyber_zeta[224], kyber_zeta[112]};
assign kyber_ntt_twiddle_mem[70] = {kyber_zeta[227], kyber_zeta[226], kyber_zeta[113]};
assign kyber_ntt_twiddle_mem[71] = {kyber_zeta[229], kyber_zeta[228], kyber_zeta[114]};
assign kyber_ntt_twiddle_mem[72] = {kyber_zeta[231], kyber_zeta[230], kyber_zeta[115]};
assign kyber_ntt_twiddle_mem[73] = {kyber_zeta[233], kyber_zeta[232], kyber_zeta[116]};
assign kyber_ntt_twiddle_mem[74] = {kyber_zeta[235], kyber_zeta[234], kyber_zeta[117]};
assign kyber_ntt_twiddle_mem[75] = {kyber_zeta[237], kyber_zeta[236], kyber_zeta[118]};
assign kyber_ntt_twiddle_mem[76] = {kyber_zeta[239], kyber_zeta[238], kyber_zeta[119]};
assign kyber_ntt_twiddle_mem[77] = {kyber_zeta[241], kyber_zeta[240], kyber_zeta[120]};
assign kyber_ntt_twiddle_mem[78] = {kyber_zeta[243], kyber_zeta[242], kyber_zeta[121]};
assign kyber_ntt_twiddle_mem[79] = {kyber_zeta[245], kyber_zeta[244], kyber_zeta[122]};
assign kyber_ntt_twiddle_mem[80] = {kyber_zeta[247], kyber_zeta[246], kyber_zeta[123]};
assign kyber_ntt_twiddle_mem[81] = {kyber_zeta[249], kyber_zeta[248], kyber_zeta[124]};
assign kyber_ntt_twiddle_mem[82] = {kyber_zeta[251], kyber_zeta[250], kyber_zeta[125]};
assign kyber_ntt_twiddle_mem[83] = {kyber_zeta[253], kyber_zeta[252], kyber_zeta[126]};
assign kyber_ntt_twiddle_mem[84] = {kyber_zeta[255], kyber_zeta[254], kyber_zeta[127]};
//--------------------------------------------------------

assign kyber_intt_twiddle_mem[0]  = {kyber_zetainv[127], kyber_zetainv[254], kyber_zetainv[255]};
assign kyber_intt_twiddle_mem[1]  = {kyber_zetainv[126], kyber_zetainv[252], kyber_zetainv[253]};
assign kyber_intt_twiddle_mem[2]  = {kyber_zetainv[125], kyber_zetainv[250], kyber_zetainv[251]};
assign kyber_intt_twiddle_mem[3]  = {kyber_zetainv[124], kyber_zetainv[248], kyber_zetainv[249]};
assign kyber_intt_twiddle_mem[4]  = {kyber_zetainv[123], kyber_zetainv[246], kyber_zetainv[247]};
assign kyber_intt_twiddle_mem[5]  = {kyber_zetainv[122], kyber_zetainv[244], kyber_zetainv[245]};
assign kyber_intt_twiddle_mem[6]  = {kyber_zetainv[121], kyber_zetainv[242], kyber_zetainv[243]};
assign kyber_intt_twiddle_mem[7]  = {kyber_zetainv[120], kyber_zetainv[240], kyber_zetainv[241]};
assign kyber_intt_twiddle_mem[8]  = {kyber_zetainv[119], kyber_zetainv[238], kyber_zetainv[239]};
assign kyber_intt_twiddle_mem[9]  = {kyber_zetainv[118], kyber_zetainv[236], kyber_zetainv[237]};
assign kyber_intt_twiddle_mem[10] = {kyber_zetainv[117], kyber_zetainv[234], kyber_zetainv[235]};
assign kyber_intt_twiddle_mem[11] = {kyber_zetainv[116], kyber_zetainv[232], kyber_zetainv[233]};
assign kyber_intt_twiddle_mem[12] = {kyber_zetainv[115], kyber_zetainv[230], kyber_zetainv[231]};
assign kyber_intt_twiddle_mem[13] = {kyber_zetainv[114], kyber_zetainv[228], kyber_zetainv[229]};
assign kyber_intt_twiddle_mem[14] = {kyber_zetainv[113], kyber_zetainv[226], kyber_zetainv[227]};
assign kyber_intt_twiddle_mem[15] = {kyber_zetainv[112], kyber_zetainv[224], kyber_zetainv[225]};
assign kyber_intt_twiddle_mem[16] = {kyber_zetainv[111], kyber_zetainv[222], kyber_zetainv[223]};
assign kyber_intt_twiddle_mem[17] = {kyber_zetainv[110], kyber_zetainv[220], kyber_zetainv[221]};
assign kyber_intt_twiddle_mem[18] = {kyber_zetainv[109], kyber_zetainv[218], kyber_zetainv[219]};
assign kyber_intt_twiddle_mem[19] = {kyber_zetainv[108], kyber_zetainv[216], kyber_zetainv[217]};
assign kyber_intt_twiddle_mem[20] = {kyber_zetainv[107], kyber_zetainv[214], kyber_zetainv[215]};
assign kyber_intt_twiddle_mem[21] = {kyber_zetainv[106], kyber_zetainv[212], kyber_zetainv[213]};
assign kyber_intt_twiddle_mem[22] = {kyber_zetainv[105], kyber_zetainv[210], kyber_zetainv[211]};
assign kyber_intt_twiddle_mem[23] = {kyber_zetainv[104], kyber_zetainv[208], kyber_zetainv[209]};
assign kyber_intt_twiddle_mem[24] = {kyber_zetainv[103], kyber_zetainv[206], kyber_zetainv[207]};
assign kyber_intt_twiddle_mem[25] = {kyber_zetainv[102], kyber_zetainv[204], kyber_zetainv[205]};
assign kyber_intt_twiddle_mem[26] = {kyber_zetainv[101], kyber_zetainv[202], kyber_zetainv[203]};
assign kyber_intt_twiddle_mem[27] = {kyber_zetainv[100], kyber_zetainv[200], kyber_zetainv[201]};
assign kyber_intt_twiddle_mem[28] = {kyber_zetainv[99], kyber_zetainv[198], kyber_zetainv[199]};
assign kyber_intt_twiddle_mem[29] = {kyber_zetainv[98], kyber_zetainv[196], kyber_zetainv[197]};
assign kyber_intt_twiddle_mem[30] = {kyber_zetainv[97], kyber_zetainv[194], kyber_zetainv[195]};
assign kyber_intt_twiddle_mem[31] = {kyber_zetainv[96], kyber_zetainv[192], kyber_zetainv[193]};
assign kyber_intt_twiddle_mem[32] = {kyber_zetainv[95], kyber_zetainv[190], kyber_zetainv[191]};
assign kyber_intt_twiddle_mem[33] = {kyber_zetainv[94], kyber_zetainv[188], kyber_zetainv[189]};
assign kyber_intt_twiddle_mem[34] = {kyber_zetainv[93], kyber_zetainv[186], kyber_zetainv[187]};
assign kyber_intt_twiddle_mem[35] = {kyber_zetainv[92], kyber_zetainv[184], kyber_zetainv[185]};
assign kyber_intt_twiddle_mem[36] = {kyber_zetainv[91], kyber_zetainv[182], kyber_zetainv[183]};
assign kyber_intt_twiddle_mem[37] = {kyber_zetainv[90], kyber_zetainv[180], kyber_zetainv[181]};
assign kyber_intt_twiddle_mem[38] = {kyber_zetainv[89], kyber_zetainv[178], kyber_zetainv[179]};
assign kyber_intt_twiddle_mem[39] = {kyber_zetainv[88], kyber_zetainv[176], kyber_zetainv[177]};
assign kyber_intt_twiddle_mem[40] = {kyber_zetainv[87], kyber_zetainv[174], kyber_zetainv[175]};
assign kyber_intt_twiddle_mem[41] = {kyber_zetainv[86], kyber_zetainv[172], kyber_zetainv[173]};
assign kyber_intt_twiddle_mem[42] = {kyber_zetainv[85], kyber_zetainv[170], kyber_zetainv[171]};
assign kyber_intt_twiddle_mem[43] = {kyber_zetainv[84], kyber_zetainv[168], kyber_zetainv[169]};
assign kyber_intt_twiddle_mem[44] = {kyber_zetainv[83], kyber_zetainv[166], kyber_zetainv[167]};
assign kyber_intt_twiddle_mem[45] = {kyber_zetainv[82], kyber_zetainv[164], kyber_zetainv[165]};
assign kyber_intt_twiddle_mem[46] = {kyber_zetainv[81], kyber_zetainv[162], kyber_zetainv[163]};
assign kyber_intt_twiddle_mem[47] = {kyber_zetainv[80], kyber_zetainv[160], kyber_zetainv[161]};
assign kyber_intt_twiddle_mem[48] = {kyber_zetainv[79], kyber_zetainv[158], kyber_zetainv[159]};
assign kyber_intt_twiddle_mem[49] = {kyber_zetainv[78], kyber_zetainv[156], kyber_zetainv[157]};
assign kyber_intt_twiddle_mem[50] = {kyber_zetainv[77], kyber_zetainv[154], kyber_zetainv[155]};
assign kyber_intt_twiddle_mem[51] = {kyber_zetainv[76], kyber_zetainv[152], kyber_zetainv[153]};
assign kyber_intt_twiddle_mem[52] = {kyber_zetainv[75], kyber_zetainv[150], kyber_zetainv[151]};
assign kyber_intt_twiddle_mem[53] = {kyber_zetainv[74], kyber_zetainv[148], kyber_zetainv[149]};
assign kyber_intt_twiddle_mem[54] = {kyber_zetainv[73], kyber_zetainv[146], kyber_zetainv[147]};
assign kyber_intt_twiddle_mem[55] = {kyber_zetainv[72], kyber_zetainv[144], kyber_zetainv[145]};
assign kyber_intt_twiddle_mem[56] = {kyber_zetainv[71], kyber_zetainv[142], kyber_zetainv[143]};
assign kyber_intt_twiddle_mem[57] = {kyber_zetainv[70], kyber_zetainv[140], kyber_zetainv[141]};
assign kyber_intt_twiddle_mem[58] = {kyber_zetainv[69], kyber_zetainv[138], kyber_zetainv[139]};
assign kyber_intt_twiddle_mem[59] = {kyber_zetainv[68], kyber_zetainv[136], kyber_zetainv[137]};
assign kyber_intt_twiddle_mem[60] = {kyber_zetainv[67], kyber_zetainv[134], kyber_zetainv[135]};
assign kyber_intt_twiddle_mem[61] = {kyber_zetainv[66], kyber_zetainv[132], kyber_zetainv[133]};
assign kyber_intt_twiddle_mem[62] = {kyber_zetainv[65], kyber_zetainv[130], kyber_zetainv[131]};
assign kyber_intt_twiddle_mem[63] = {kyber_zetainv[64], kyber_zetainv[128], kyber_zetainv[129]};
assign kyber_intt_twiddle_mem[64] = {kyber_zetainv[31], kyber_zetainv[62], kyber_zetainv[63]};
assign kyber_intt_twiddle_mem[65] = {kyber_zetainv[30], kyber_zetainv[60], kyber_zetainv[61]};
assign kyber_intt_twiddle_mem[66] = {kyber_zetainv[29], kyber_zetainv[58], kyber_zetainv[59]}; 
assign kyber_intt_twiddle_mem[67] = {kyber_zetainv[28], kyber_zetainv[56], kyber_zetainv[57]};
assign kyber_intt_twiddle_mem[68] = {kyber_zetainv[27], kyber_zetainv[54], kyber_zetainv[55]};
assign kyber_intt_twiddle_mem[69] = {kyber_zetainv[26], kyber_zetainv[52], kyber_zetainv[53]};
assign kyber_intt_twiddle_mem[70] = {kyber_zetainv[25], kyber_zetainv[50], kyber_zetainv[51]};
assign kyber_intt_twiddle_mem[71] = {kyber_zetainv[24], kyber_zetainv[48], kyber_zetainv[49]};
assign kyber_intt_twiddle_mem[72] = {kyber_zetainv[23], kyber_zetainv[46], kyber_zetainv[47]};
assign kyber_intt_twiddle_mem[73] = {kyber_zetainv[22], kyber_zetainv[44], kyber_zetainv[45]};
assign kyber_intt_twiddle_mem[74] = {kyber_zetainv[21], kyber_zetainv[42], kyber_zetainv[43]};
assign kyber_intt_twiddle_mem[75] = {kyber_zetainv[20], kyber_zetainv[40], kyber_zetainv[41]};
assign kyber_intt_twiddle_mem[76] = {kyber_zetainv[19], kyber_zetainv[38], kyber_zetainv[39]};
assign kyber_intt_twiddle_mem[77] = {kyber_zetainv[18], kyber_zetainv[36], kyber_zetainv[37]};
assign kyber_intt_twiddle_mem[78] = {kyber_zetainv[17], kyber_zetainv[34], kyber_zetainv[35]};
assign kyber_intt_twiddle_mem[79] = {kyber_zetainv[16], kyber_zetainv[32], kyber_zetainv[33]};
assign kyber_intt_twiddle_mem[80] = {kyber_zetainv[7], kyber_zetainv[14], kyber_zetainv[15]};
assign kyber_intt_twiddle_mem[81] = {kyber_zetainv[6], kyber_zetainv[12], kyber_zetainv[13]};
assign kyber_intt_twiddle_mem[82] = {kyber_zetainv[5], kyber_zetainv[10], kyber_zetainv[11]};
assign kyber_intt_twiddle_mem[83] = {kyber_zetainv[4], kyber_zetainv[8], kyber_zetainv[9]};
assign kyber_intt_twiddle_mem[84] = {kyber_zetainv[1], kyber_zetainv[2], kyber_zetainv[3]};

endmodule