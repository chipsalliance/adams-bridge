// `include "$COMPILE_ROOT/utb/sequences/ntt_seq/ntt_base_seq.sv"
// `include "$COMPILE_ROOT/utb/sequences/ntt_seq/ntt_fwd_seq.sv"
