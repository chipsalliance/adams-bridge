// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
//======================================================================
//
// Module: abr_masked_A2B_conv
// Description: This module implements a pipelined, parametric ripple-carry adder using the abr_masked_full_adder.
//              It performs addition of two boolean shared inputs, producing a boolean shared output.
// 
// Parameters:
//  - WIDTH: Specifies the bit-width of the operands.
// 
// Functionality:
//  - The module performs a share conversion between arithmetic and Boolean shares.
//  - It takes WIDTH+2 cycle latency
//
//======================================================================

 module abr_masked_A2B_conv #(
    parameter WIDTH = 8 // Default width is 8 bits
)(
    input wire clk,                                 // Clock signal
    input wire rst_n,                               // Active low reset signal
    input wire zeroize,                             // Zeroize signal
    input wire [1:0] x [WIDTH-1:0],                 // WIDTH-bit arithmetic shares operand x
    input wire [WIDTH-1:0] rnd,                     // Random bits for masking
    input wire [WIDTH-1:0] rnd_for_Boolean0,        // Random bits for masking
    input wire [WIDTH-1:0] rnd_for_Boolean1,        // Random bits for masking

    output logic [1:0] s [WIDTH-1:0]
);

    // Internal signals
    logic [1:0] carry [WIDTH:0]; // Carry signals for each stage
    logic [1:0] sum [WIDTH-1:0]; // Sum signals for each stage
    logic [1:0] x_reg [WIDTH-1:0][WIDTH-1:0]; // Pipeline registers for x
    logic [1:0] y_reg [WIDTH-1:0][WIDTH-1:0]; // Pipeline registers for y
    logic [1:0] sum_reg [WIDTH-1:0][WIDTH-1:0]; // Pipeline registers for sum
    logic [1:0] the_last_sum;

    // Initialize the first carry input to 0
    assign carry[0] = 2'b00;

    // Generate the full adders for each bit
    genvar i;
    generate
        for (i = 0; i < WIDTH; i = i + 1) begin : gen_full_adders
            // Pipeline registers for x and y inputs
            always_ff @(posedge clk or negedge rst_n) begin
                if (!rst_n) begin
                    for (int j = 0; j < WIDTH; j = j + 1) begin
                        x_reg[i][j] <= 2'b00;
                        y_reg[i][j] <= 2'b00;
                    end
                end
                else if (zeroize) begin
                    for (int j = 0; j < WIDTH; j = j + 1) begin
                        x_reg[i][j] <= 2'b00;
                        y_reg[i][j] <= 2'b00;
                    end
                end
                else begin
                    for (int j = 0; j < WIDTH; j = j + 1) begin
                        if (j == 0) begin
                            x_reg[i][j] <= {rnd_for_Boolean0[i], (x[i][0] ^ rnd_for_Boolean0[i])};
                            y_reg[i][j] <= {rnd_for_Boolean1[i], (x[i][1] ^ rnd_for_Boolean1[i])};
                        end
                        else begin
                            x_reg[i][j] <= x_reg[i][j-1];
                            y_reg[i][j] <= y_reg[i][j-1];
                        end
                    end
                end
            end

            // Pipeline registers for sum output
            always_ff @(posedge clk or negedge rst_n) begin
                if (!rst_n) begin
                    for (int j = 0; j < WIDTH; j = j + 1) begin
                        sum_reg[i][j] <= 2'b00;
                    end
                end
                else if (zeroize) begin
                    for (int j = 0; j < WIDTH; j = j + 1) begin
                        sum_reg[i][j] <= 2'b00;
                    end
                end
                else begin
                    for (int j = i; j < WIDTH; j = j + 1) begin
                        if (j == i && i == WIDTH-1) begin
                            sum_reg[i][j] <= the_last_sum;
                        end
                        else if (j == i) begin
                            sum_reg[i][j] <= sum[i];
                        end
                        else begin
                            sum_reg[i][j] <= sum_reg[i][j-1];
                        end
                    end
                end
            end
            if (i<(WIDTH-1)) begin
                // Instance of abr_masked_full_adder
                abr_masked_full_adder u_abr_masked_full_adder (
                    .clk(clk),              // Connect clk to clk
                    .rst_n(rst_n),          // Connect rst_n to rst_n
                    .zeroize(zeroize),      // Connect zeroize to zeroize
                    .x(x_reg[i][i]),  // Connect x to the last stage of the x pipeline
                    .y(y_reg[i][i]),  // Connect y to the last stage of the y pipeline
                    .c_in(carry[i]),        // Connect c_in to carry[i]
                    .rnd(rnd[i]),           // Connect rnd to corresponding random bit
                    .s(sum[i]),             // Connect sum to sum[i]
                    .c_out(carry[i+1])      // Connect carry out to carry[i+1]
                );
            end
        end
    endgenerate

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            the_last_sum    <= 2'b00;
        end
        else if (zeroize) begin
            the_last_sum    <= 2'b00;
        end
        else begin
            the_last_sum <= x_reg[WIDTH-1][WIDTH-1] ^ y_reg[WIDTH-1][WIDTH-1] ^ carry[WIDTH-1];
        end
    end

    // Assign the outputs
    always_comb begin
        for (int i =0; i<WIDTH; i++) begin
            s[i] = sum_reg[i][WIDTH-1];
        end
    end

endmodule : abr_masked_A2B_conv
