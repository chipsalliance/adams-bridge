//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This file contains the top level sequence used in  example_derived_test.
// It is an example of a sequence that is extended from %(benchName)_bench_sequence_base
// and can override %(benchName)_bench_sequence_base.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

typedef struct {
  string seed_d;       // Input SEED_D
  string seed_z;       // Input SEED_Z
  string expected_PK;  // Expected Public Key
  string expected_SK;  // Expected Secret Key
} mlkem_keygen_kat_t;

class ML_KEM_keygen_KATs_sequence extends mldsa_bench_sequence_base;

  `uvm_object_utils(ML_KEM_keygen_KATs_sequence);

    
    // KAT arrays
  mlkem_keygen_kat_t keygen_kats[];
  bit [31:0] kat_seed_d [];
  bit [31:0] kat_seed_z [];
  bit ready;
  bit valid;
  int value;
  

  function new(string name = "");
    super.new(name);
    keygen_kats = new[1];
    kat_seed_d = new[8];
    kat_seed_z = new[8];
  endfunction

  virtual task body();
    reg_model.reset();
    #400;


    if (reg_model.default_map == null) begin
      `uvm_fatal("MAP_ERROR", "mldsa_uvm_rm.default_map map is not initialized");
    end else begin
      `uvm_info("MAP_INIT", "mldsa_uvm_rm.default_map is initialized", UVM_LOW);
    end

    
   // KeyGen KATs
    keygen_kats[0].seed_d = "CDF4E658BDD4636F09F70BD76CE6D1AF028562586EF237C7481033EE03C31FF2";
    keygen_kats[0].seed_z = "38CD80FE6CD34678DE86E55E145BAF191B675C19C485C54EF3522C044D42F6EE";
    keygen_kats[0].expected_PK = "B1B5987867073BA270695AB4FC076975CC5C1BE18F8DCC36660ACE35A72D678639483C86B780A483FB3C77C8998F7047CC027CE6522998D796E8F288EA893D3E34ACB1CB4375657819012BAADB7B8A878F8FD4C7B6B42641F5B1C286ACBB41783B2CBE62A167F92A274A4763A2C293360179421CCC933B96A8C693FE47730DB1450FE04DC98B8C4E05B6A10B5CF07B44A620C3576932BA420BC536C149D1BA3CB40DF2497A7E9CC8E385A291C411717368180AA4AA00026C08B1A051A0B0C6BA96572AF9511FF020A32F47CB2EA4A9428345AC347CE1968A1159847F2B2D46355C63FB5043765F37E967A97B2113E52A66C3C8D1F3127814553516BFA2BCB26B537F1FD23CFAEAC28D842CF334534FE24782D7841BC3C0E2A9721D7084FAA32F03B00F018028A9F650136C79E6A39DCEF08D23B1B936A2A2B5790022EB8184052A2D39898761289F13BC587898F4538ACA0B19C471BB7DCA949A478FE7D36A71A8BAB72976EABA62BAFAB2BF772EE48CC12B63C06BE90929E562925562803903A4C1CAE1984A82D95A3A507608C337A3F7B89FC09883DA24B8E3ABB3789D1CA938C0E747FA1A38153B96D1122DC6B69258F474324A3A7024713B9CC896118F09087B52BC079277B0B9004B45330707AC5E1E8C34CBC40971D8ACC49C93A5903A9394CA873A7E7AF09CE2192BEC9A6070D28118715B5EC592481BBDDB67C14ACB88823B7161E85798A36AD7B68AE5584FA02C66EE7A6A35A97D496C8E9927421B110E00468729D5924D016A68800CCCA3AEDE4CCC6471C07C2A0B8B5168B4647CB240AC8745C22B0AADE8B4883A7A43F53ABE21B384BA94741A787634E72B599C25D3904627C69B91013A4AE749117B0F41AA86B389BF46707D07812B7424B3E5F1BA000C9D1386091C29337AD697E3089D2D5146FD1BBF66ECCAE1430EEC8A1308CB99210C19A71B3A0DF42559C4A7EC7BA901C3BB6168B5CCE02989E54DC193229759B9FE3B5E31013117DCB67EE53201E18F52931239B7A2FD477970CBA3D0621CD555C498600759746453C94FBC539608F4B47631B3A6C4AB32849F8716A557B93A417DB8FBC47945B60765D6D59FCED9312E8435B43711118891E6EEB2C1";
    keygen_kats[0].expected_SK = "6441B2F8804D0D9B08827A6E8AA3B25032BA71E341297BBAA3F33835149825D2810182C9A24B0892355F68CC3719B2085CD2B205910F450A0D4F4CB49AC0A826B88BBDBAC1429C6AF3E25E67338D3525658E5433A7CBA2CAC6CC07933A3BB1BBD7A10E87B481EA54A43EC926B82044FAC0895C1B3535669C77139729763CBE466BCCFCA940AC3734070B88B7C3D944B3D465188644819A9A8A413C9D8911668C4B567EAC80531CADC8717549C483BB39866EB68EB8E2AE53836D893864B7CCBE519893C8F7CAC00B2AE30C059E54A09799273DF44F2C8CBD426C618BDB676CC26073D46D9E652EE6A667A5F0CD60E54E9D22CFC2A2CA23D39040A38873646293CCAF2BB9110DD217B0EB065E7737A4B85CA6A73C215C0D2B899B01B30E461009E28CA280AB6805FC2A91C6CB665194D7430640F65A87714BB8632718B94EA649A95BB80DAD67134BB8628A6790C5E9013939306D8649AA65B67260BD6D28BE682562352935A95839AD672059D9C30794C513A5726EDB962E385A71A76A9454BBDB9C2E45315C3D07298C19015D68347D7067582B3B8F8CB59AE582AE4B2C74AC6AD894330F93B18571976E01AD9DE592CAFAC2805712AEB60351989946C13F831327AA120C8A368BBFBA7A8999B3B9E762E700227E0B4D0E7C00603768FA237068D95B5B0045BC1206381B5E9175460F31855FB4BF2C2376C0E515A6224D3BF94A099A89FC215F9C39958C440FF8EB71A4476C9C4C4357045547182A537181ED48B07C275170C853C08C71CD5C2E526700688C394E166062EC35A5B062A31306BB5C30224BCA7E1664DCD3C1061141CFE83714449FEFCA2A792B734AC247CA3479C0A469F763AABAA6331D413201699B2AE22A79F076C6F2C1BEE8AFF3D3960CC37A242391484C8FF872C65D576E05CA0E7F614A3DD43D8E23658699960773178BE97F2E96BE4DA5530C3A7DEC06346A092860458681024969A16A3CF128D4439DF9780F38F16F89848299416A0C5460600A517D615DCDA4204D36C167BB083272C69977A175F3B434DB79724A6C51279428CA6BB8476CCC2C23033C768B1628B1B5987867073BA270695AB4FC076975CC5C1BE18F8DCC36660ACE35A72D678639483C86B780A483FB3C77C8998F7047CC027CE6522998D796E8F288EA893D3E34ACB1CB4375657819012BAADB7B8A878F8FD4C7B6B42641F5B1C286ACBB41783B2CBE62A167F92A274A4763A2C293360179421CCC933B96A8C693FE47730DB1450FE04DC98B8C4E05B6A10B5CF07B44A620C3576932BA420BC536C149D1BA3CB40DF2497A7E9CC8E385A291C411717368180AA4AA00026C08B1A051A0B0C6BA96572AF9511FF020A32F47CB2EA4A9428345AC347CE1968A1159847F2B2D46355C63FB5043765F37E967A97B2113E52A66C3C8D1F3127814553516BFA2BCB26B537F1FD23CFAEAC28D842CF334534FE24782D7841BC3C0E2A9721D7084FAA32F03B00F018028A9F650136C79E6A39DCEF08D23B1B936A2A2B5790022EB8184052A2D39898761289F13BC587898F4538ACA0B19C471BB7DCA949A478FE7D36A71A8BAB72976EABA62BAFAB2BF772EE48CC12B63C06BE90929E562925562803903A4C1CAE1984A82D95A3A507608C337A3F7B89FC09883DA24B8E3ABB3789D1CA938C0E747FA1A38153B96D1122DC6B69258F474324A3A7024713B9CC896118F09087B52BC079277B0B9004B45330707AC5E1E8C34CBC40971D8ACC49C93A5903A9394CA873A7E7AF09CE2192BEC9A6070D28118715B5EC592481BBDDB67C14ACB88823B7161E85798A36AD7B68AE5584FA02C66EE7A6A35A97D496C8E9927421B110E00468729D5924D016A68800CCCA3AEDE4CCC6471C07C2A0B8B5168B4647CB240AC8745C22B0AADE8B4883A7A43F53ABE21B384BA94741A787634E72B599C25D3904627C69B91013A4AE749117B0F41AA86B389BF46707D07812B7424B3E5F1BA000C9D1386091C29337AD697E3089D2D5146FD1BBF66ECCAE1430EEC8A1308CB99210C19A71B3A0DF42559C4A7EC7BA901C3BB6168B5CCE02989E54DC193229759B9FE3B5E31013117DCB67EE53201E18F52931239B7A2FD477970CBA3D0621CD555C498600759746453C94FBC539608F4B47631B3A6C4AB32849F8716A557B93A417DB8FBC47945B60765D6D59FCED9312E8435B43711118891E6EEB2C173EAB9578A8556AA31C7CDC35F49987E3F6E1843CA41137BF1D50DC20557F4DF38CD80FE6CD34678DE86E55E145BAF191B675C19C485C54EF3522C044D42F6EE";

    // Iterate through KATs and validate
    foreach (keygen_kats[i]) begin
      parse_hex_to_array(keygen_kats[i].seed_d, kat_seed_d);
      parse_hex_to_array(keygen_kats[i].seed_z, kat_seed_z);
      parse_hex_to_array(keygen_kats[i].expected_PK, PK);
      parse_hex_to_array(keygen_kats[i].expected_SK, SK);

      `uvm_info("KAT", $sformatf("Running KeyGen KAT %0d", i), UVM_LOW);

      // Wait for ready flag in MLKEM_STATUS
      ready = 0;
      while (!ready) begin
        reg_model.MLKEM_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ_FAIL", "Failed to read MLKEM_STATUS");
        end else begin
          `uvm_info("REG_READ_PASS", $sformatf("MLKEM_STATUS: %h", data), UVM_HIGH);
        end
        ready = data[0];
      end

      // Write SEED to ML_KEM_SEED_D registers
      foreach (reg_model.MLKEM_SEED_D[j]) begin
        reg_model.MLKEM_SEED_D[j].write(status, kat_seed_d[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLKEM_SEED_D[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLKEM_SEED_D[%0d]: %h", j, kat_seed_d[j]), UVM_LOW);
        end
      end

      // Write SEED to ML_KEM_SEED_Z registers
      foreach (reg_model.MLKEM_SEED_Z[j]) begin
        reg_model.MLKEM_SEED_Z[j].write(status, kat_seed_z[j], UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_WRITE_FAIL", $sformatf("Failed to write MLKEM_SEED_Z[%0d] for KAT %0d", j, i));
        end else begin
          `uvm_info("REG_WRITE_PASS", $sformatf("Successfully wrote MLKEM_SEED_Z[%0d]: %h", j, kat_seed_z[j]), UVM_LOW);
        end
      end

      // Trigger KeyGen operation
      data = 'h00000001; // KeyGen command
      reg_model.MLKEM_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE_FAIL", "Failed to write MLKEM_CTRL to trigger KeyGen");
      end else begin
        `uvm_info("REG_WRITE_PASS", "Successfully wrote MLKEM_CTRL to trigger KeyGen", UVM_LOW);
      end

      // Wait for ready flag in MLKEM_STATUS
      valid =0;
      while(!valid) begin
        reg_model.MLKEM_STATUS.read(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_STATUS"));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_STATUS: %0h", data), UVM_HIGH);
        end
        valid = data[1];
      end

      // Reading MLKEM_ENCAPS_KEY register
      for(int i = 0; i < reg_model.MLKEM_ENCAPS_KEY.m_mem.get_size(); i++) begin
        reg_model.MLKEM_ENCAPS_KEY.m_mem.read(status, i, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_ENCAPS_KEY[%0d]", i));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_ENCAPS_KEY[%0d]: %0h", i, data), UVM_LOW);
          if (PK[i] != data)
          `uvm_error("REG_READ", $sformatf("MLKEM_ENCAPS_KEY[%0d] mismatch: actual=0x%08h, expected=0x%08h",
                    i, data, PK[i]));
        end
      end

      // Reading MLKEM_DECAPS_KEY register
      for(int i = 0; i < reg_model.MLKEM_DECAPS_KEY.m_mem.get_size(); i++) begin
        reg_model.MLKEM_DECAPS_KEY.m_mem.read(status, i, data, UVM_FRONTDOOR, reg_model.default_map, this);
        if (status != UVM_IS_OK) begin
          `uvm_error("REG_READ", $sformatf("Failed to read MLKEM_DECAPS_KEY[%0d]", i));
        end else begin
          `uvm_info("REG_READ", $sformatf("MLKEM_DECAPS_KEY[%0d]: %0h", i, data), UVM_LOW);
          if (SK[i] != data)
          `uvm_error("REG_READ", $sformatf("MLKEM_DECAPS_KEY[%0d] mismatch: actual=0x%08h, expected=0x%08h",
                    i, data, SK[i]));
        end
      end

      data = 'h0000_0008; // Perform zeorization operation
      reg_model.MLDSA_CTRL.write(status, data, UVM_FRONTDOOR, reg_model.default_map, this);
      if (status != UVM_IS_OK) begin
        `uvm_error("REG_WRITE", $sformatf("Failed to write MLDSA_CTRL"));
      end else begin
        `uvm_info("REG_WRITE", $sformatf("MLDSA_CTRL written with %0h and zeroized", data), UVM_LOW);
      end
    end

    `uvm_info("KAT", $sformatf("KeyGen KAT validation completed"), UVM_LOW);


  endtask

   


  endclass




// pragma uvmf custom external begin
// pragma uvmf custom external end



